module sprite_tile(
	output logic [23:0] mem [0:4899],
	output logic [23:0] mem_red [0:4899],
	output logic [23:0] mem_yellow [0:4899],
	output logic [23:0] mem_green [0:4899]
	);

logic [23:0] memory [0:4899] = '{
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011011010001,
    24'b000000010110011011010001,
    24'b000000010110011011010000,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011001111,
    24'b000000000110011011001111,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010001,
    24'b000000010110011011010001,
    24'b000000010110011011010001,
    24'b000000010110011011010001,
    24'b000000010110011011010001,
    24'b000000000110100011001110,
    24'b000000000110100011001110,
    24'b000000000110011111001110,
    24'b000000010110100011001101,
    24'b000000000110011111001110,
    24'b000000000110011111001101,
    24'b000000000110011111001100,
    24'b000000010110011111001100,
    24'b000000010110011111001100,
    24'b000000000110011111001100,
    24'b000000000110100011001100,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000100110011111001111,
    24'b000000100110011111001111,
    24'b000000100110011111010001,
    24'b000000010110011011010000,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000000110100011010011,
    24'b000000000110100011010011,
    24'b000000000110100011010001,
    24'b000000000110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000010110100011010001,
    24'b000000010110100011001111,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000010110011011001111,
    24'b000000010110011011001111,
    24'b000000100110011011001110,
    24'b000000010110011011001111,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111001110,
    24'b000000100110100011001110,
    24'b000000010110011011001111,
    24'b000000100110011111010010,
    24'b000000100110011011010100,
    24'b000000100110011011010101,
    24'b000000000110011111010011,
    24'b000000000110100011010010,
    24'b000000010110011111010001,
    24'b000000010110011111010000,
    24'b000000110110011111001111,
    24'b000000100110011111001111,
    24'b000000010110011111001111,
    24'b000000010110011111001100,
    24'b000000010110011111001100,
    24'b000000100110100111001110,
    24'b000000110110100111010010,
    24'b000001000110100111010100,
    24'b000000100110011111010010,
    24'b000000100110100011010100,
    24'b000000010110011111010011,
    24'b000000100110011111010100,
    24'b000000100110011111010100,
    24'b000000100110011111010011,
    24'b000001000110011011010011,
    24'b000001000110011011010011,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111001100,
    24'b000000000110011011001011,
    24'b000000010110011011001110,
    24'b000000010110011011010010,
    24'b000000010110010111010100,
    24'b000000000110010011010100,
    24'b000000010110100011010001,
    24'b000000010110011011001111,
    24'b000001000110011111001111,
    24'b000001000110011011001100,
    24'b000001000110010111001011,
    24'b000001000110010111001011,
    24'b000001010110011011001011,
    24'b000001000110010111000110,
    24'b000001000110010111000101,
    24'b000001010110011011001000,
    24'b000001010110010111001011,
    24'b000001000110010111001011,
    24'b000001000110011011001011,
    24'b000000110110011011001101,
    24'b000001000110011011010000,
    24'b000000110110010111010000,
    24'b000000010110011011010001,
    24'b000000110110011011010000,
    24'b000001000110011011010001,
    24'b000001000110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000100110011111010000,
    24'b000000010110011011001110,
    24'b000000000110010111001110,
    24'b000000010110011111010001,
    24'b000001000110101111010111,
    24'b000000110110100111010100,
    24'b000000100110010011001100,
    24'b000001000110011011001011,
    24'b000001110110011011000111,
    24'b000010110110001111000001,
    24'b000100100110001111000000,
    24'b000100110110001010111100,
    24'b000100000101111010110110,
    24'b000100010101101110110011,
    24'b000100000101101110101111,
    24'b000100000101101110101101,
    24'b000100000101101110101111,
    24'b000101000101111010110111,
    24'b000011110110010110111100,
    24'b000010010110001010111010,
    24'b000010010110010011000001,
    24'b000001100110010111000101,
    24'b000001000110010011001010,
    24'b000001010110010111001111,
    24'b000001000110011111001011,
    24'b000001000110011111001111,
    24'b000000110110100011010001,
    24'b000000010110011011001111,
    24'b000000000110011111001111,
    24'b000000000110100011010001,
    24'b000000000110011111010000,
    24'b000000100110011011001110,
    24'b000000000110100011010010,
    24'b000000000110100011010010,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110100011010010,
    24'b000000000110011111001111,
    24'b000000110110010111001010,
    24'b000000000110010111001111,
    24'b000000110110100111010001,
    24'b000001000110010011001001,
    24'b000011000110100011001011,
    24'b000001110110000111000100,
    24'b000100010110011011000110,
    24'b000101010110001110111011,
    24'b001000100101011110011100,
    24'b000100010011111001111000,
    24'b000001110010011101010110,
    24'b000000000001011100111010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001000000110011,
    24'b000000000001110101001001,
    24'b000010010011010101101000,
    24'b000101000100111110001100,
    24'b000101110101111010101001,
    24'b000100110110000110111010,
    24'b000011110110001111001001,
    24'b000001000110010111001100,
    24'b000000100110100111001111,
    24'b000001000110101011010000,
    24'b000000010110011011010000,
    24'b000000000110011011010100,
    24'b000000000110011111001111,
    24'b000000000110100011001011,
    24'b000000000110100011010001,
    24'b000000000110011011010010,
    24'b000000110110011011001100,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000000110011011010010,
    24'b000000110110011011001101,
    24'b000001010110011011001101,
    24'b000000000110100011010100,
    24'b000000000110100011010101,
    24'b000010110110010111001000,
    24'b000111110110000010110000,
    24'b001000000100110110001010,
    24'b000001110010010001010011,
    24'b000000010000111100110011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000100001001100110010,
    24'b000011010011100101111000,
    24'b000111010101101110110001,
    24'b000110000110100011001100,
    24'b000010100110010011001100,
    24'b000000110110011111001001,
    24'b000000100110011011001011,
    24'b000000110110011111001010,
    24'b000000100110011011001000,
    24'b000000100110010111001100,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111001101,
    24'b000001010110100011001110,
    24'b000000000110011011010111,
    24'b000000010110101011011111,
    24'b000011010110001111000111,
    24'b000111100101110110101110,
    24'b000011110011101001111001,
    24'b000000000001000000111000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001011010010010100100011,
    24'b011101100110101101100100,
    24'b101010101001110110010101,
    24'b110100001100001110111001,
    24'b110111101101000011001000,
    24'b111001001101010111001111,
    24'b111001101101011011010000,
    24'b111001101101011011010010,
    24'b111000101101001011001111,
    24'b110111011100110011001000,
    24'b101101101011000110100110,
    24'b100011001000100010000001,
    24'b010100010100110001001010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000001000010010001010110,
    24'b000101000100111110010111,
    24'b000011010110001010111110,
    24'b000001000110101011001100,
    24'b000000110110010111001010,
    24'b000000010110001011001100,
    24'b000000000110100011010011,
    24'b000000010110110011011000,
    24'b000000010110010111010100,
    24'b000000100110010111010000,
    24'b000000100110011011010001,
    24'b000000010110011011010000,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010000,
    24'b000000000110011111001111,
    24'b000000000110011111001100,
    24'b000010000110011111001000,
    24'b000010100110011011001010,
    24'b000100010110001110111101,
    24'b000011100011111001111101,
    24'b000000010001000100101101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010100110100101101001101,
    24'b101101111010111010110000,
    24'b111000111101011011010000,
    24'b111011101101111111011001,
    24'b111100011110001011011010,
    24'b111100011110001011011001,
    24'b111100101110001011011000,
    24'b111100011110001111011000,
    24'b111011111110000111010101,
    24'b111100001110001011010110,
    24'b111100001110001011010111,
    24'b111100001110001011011000,
    24'b111100011110001111011001,
    24'b111100001110000011010110,
    24'b111100001110000011011011,
    24'b111011011110000011011101,
    24'b111011001110010111011101,
    24'b110011111100110011000011,
    24'b011110010111100001110000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000001100010010001010101,
    24'b000101000101011110100010,
    24'b000010100110100111000100,
    24'b000000100110110011010100,
    24'b000001000110010011010010,
    24'b000010100110000111001010,
    24'b000001010110011011000110,
    24'b000000110110011011001110,
    24'b000000110110011011001110,
    24'b000000010110011011010000,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000010110100011010001,
    24'b000000010110011111010001,
    24'b000001010110010111010001,
    24'b000011100110010111001001,
    24'b000101110100111010010100,
    24'b000000100001010000110010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100010100111111101111010,
    24'b110111111101010111001100,
    24'b111011101110001111011100,
    24'b111100101110001111011011,
    24'b111011001101111111010101,
    24'b111100101110010011011011,
    24'b111100011110001011011001,
    24'b111101001110010011011011,
    24'b111100011110000011010110,
    24'b111011111101110111010010,
    24'b111100011110000111010001,
    24'b111100111110000111010110,
    24'b111100111110000111010111,
    24'b111100111110001011010111,
    24'b111100111110000111010101,
    24'b111100001110000111010110,
    24'b111011101101111111011010,
    24'b111100101110001111011110,
    24'b111011111110000111011000,
    24'b111011101110000111010011,
    24'b111100011110010011010111,
    24'b111100011110001011011010,
    24'b101110111011001110101111,
    24'b010000100011110100111100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000010100011010001101001,
    24'b000101110110000010110110,
    24'b000011000110011011001111,
    24'b000001000110010111010000,
    24'b000000010110100011010010,
    24'b000001000110010111001110,
    24'b000000110110010111001110,
    24'b000000110110010111010000,
    24'b000000100110011111010001,
    24'b000000000110011111010001,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000000110010111001111,
    24'b000000000110011011010010,
    24'b000000000110011111010100,
    24'b000000010110011011001101,
    24'b000000000110011111010100,
    24'b000000000110100011010100,
    24'b000001100110100011001110,
    24'b000000110110100011010001,
    24'b000101100110001110110011,
    24'b000011100011001101101110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100001000111100001110110,
    24'b111011011101110111010101,
    24'b111101001110001111011010,
    24'b111100011110001011011000,
    24'b111100011110001011011000,
    24'b111100011110001011010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100111110000111010101,
    24'b111100101110000111010110,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100101110000111011000,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010110,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111101001110000111100001,
    24'b111101001110001111011011,
    24'b111100101110001111010110,
    24'b110001011011100110101111,
    24'b001100110010101000100111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000110001010100111011,
    24'b000110110101100010100011,
    24'b000010100110011011001011,
    24'b000001010110100011010000,
    24'b000000110110101111010100,
    24'b000000000110011011010001,
    24'b000000000110011111010010,
    24'b000001010110100011010000,
    24'b000000000110011011001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011011001110,
    24'b000000100110011111001111,
    24'b000000010110011011010000,
    24'b000000000110011011010011,
    24'b000000010110011111001101,
    24'b000000010110011011001110,
    24'b000000010110011111001100,
    24'b000000000110011111010000,
    24'b000001010110011011001001,
    24'b000110010101110010101000,
    24'b000000100010001101010100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001111010011101001000110,
    24'b111000011101011011010101,
    24'b111011011101110111010010,
    24'b111100001101111111010101,
    24'b111100111110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100011110000111011101,
    24'b111101101110001111011100,
    24'b111100011101111111010100,
    24'b111100011110001111011010,
    24'b111100001110010111011110,
    24'b100110011000111110001011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000101000101001,
    24'b000101000100010010000000,
    24'b000101010110011110111111,
    24'b000000000110101011010101,
    24'b000001010110010111001101,
    24'b000010000110010111001100,
    24'b000000110110100111001111,
    24'b000000000110011111010000,
    24'b000000010110011011001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001111,
    24'b000000010110011011010000,
    24'b000000100110011111010001,
    24'b000000110110011011001100,
    24'b000000000110011111010010,
    24'b000000010110011011001110,
    24'b000001010110000111000001,
    24'b000101000101011010011111,
    24'b000000100001011100111011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100101111000100110000100,
    24'b111010011110001011010001,
    24'b111100111110010011011101,
    24'b111100101101111011011000,
    24'b111100101110000111010111,
    24'b111100001101111111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111011111110001011010101,
    24'b111100111110001011011010,
    24'b111101001110000111011010,
    24'b111110001110011111011111,
    24'b111011001101111011010001,
    24'b111011101101110011001101,
    24'b110111001101010111001101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000011000011100101110000,
    24'b000011010110010110111111,
    24'b000011000110001011001100,
    24'b000000110110001111010001,
    24'b000000000110101111010000,
    24'b000000000110011111001110,
    24'b000000100110010111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110010111010000,
    24'b000000100110011111010000,
    24'b000000010110011111010100,
    24'b000000010110011011010100,
    24'b000001100110010011001110,
    24'b001000110101101110100011,
    24'b000000000000110100101100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110010011100000010111001,
    24'b111100101110010111011110,
    24'b111100001110010111011110,
    24'b111101001110001011011000,
    24'b111100111110000111010100,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010100,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100001110000011010001,
    24'b111011011110010011011000,
    24'b111010111110100011100001,
    24'b010010000100010101000001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000100110011101101101110,
    24'b000100110110001111000001,
    24'b000000000110100111011011,
    24'b000000100110101111010011,
    24'b000000110110011011001101,
    24'b000000010110011111010010,
    24'b000000000110011111001110,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010001,
    24'b000000000110010111010001,
    24'b000000110110100011010010,
    24'b000001000110011011001110,
    24'b000000010110011011010000,
    24'b000010100110010111000101,
    24'b000111100101111010101011,
    24'b000000010001001000110110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110101101100111011000110,
    24'b111100011110010011011110,
    24'b111010101101110011010011,
    24'b111100101110010011011001,
    24'b111011111110000111010110,
    24'b111100101110000111010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010110,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110000111010110,
    24'b111100011110001111011001,
    24'b111100001110001011011001,
    24'b111010111101111111011000,
    24'b111010101110000111100000,
    24'b011010010110010001100101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000010100011110101110010,
    24'b000011100110011010111111,
    24'b000010000110010011001111,
    24'b000001010110010111010000,
    24'b000000000110011111010011,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010011,
    24'b000000110110011111001111,
    24'b000001010110011111001110,
    24'b000001010110011111001000,
    24'b000101110110001110110001,
    24'b000000000001001100111000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110101111101000011000011,
    24'b111101001110001111010101,
    24'b111100011101110111010011,
    24'b111101001101111111010010,
    24'b111100111110001011010001,
    24'b111100011110001011011000,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000011011001,
    24'b111100111110000111010110,
    24'b111100101110001011010011,
    24'b111100101110001011010101,
    24'b111100101110000111011001,
    24'b111100011110001011011010,
    24'b111101001110001111011011,
    24'b111110011110001111011100,
    24'b111101011101111011010110,
    24'b111100001110000011011010,
    24'b011011000110010101100010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000110100100111010000100,
    24'b000011110101111111000111,
    24'b000000100110010111010011,
    24'b000000000110011111010001,
    24'b000000010110011111010101,
    24'b000000000110011011010011,
    24'b000000000110011111010001,
    24'b000000000110011111001101,
    24'b000000000110011111001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010001,
    24'b000000010110011011001110,
    24'b000000010110011011001111,
    24'b000000000110011111010100,
    24'b000010000110100011001110,
    24'b000000110110010111001011,
    24'b000100000110010111000011,
    24'b000001100010100101011110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110100001100100010111111,
    24'b111100001110001111010101,
    24'b111100001110000011010001,
    24'b111100101110001011010101,
    24'b111100011110000111010100,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110000111010111,
    24'b111100101110000011010110,
    24'b111011111101110011010101,
    24'b111100001101110011010110,
    24'b001111010011010100111000,
    24'b000000000000000000000000,
    24'b000000000000111100101001,
    24'b000110110101100110100110,
    24'b000010000110101011001000,
    24'b000001110110011011010000,
    24'b000001000110100011010110,
    24'b000000000110011011011000,
    24'b000000000110011111010001,
    24'b000000010110100011001001,
    24'b000000000110011111010000,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110100011001011,
    24'b000000010110011011001111,
    24'b000000000110001111001101,
    24'b000010100110001110111011,
    24'b000100000100001101110111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101110101010110010100101,
    24'b111100111110011011100000,
    24'b111011101101110011010011,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100011110000111010111,
    24'b111100101110000111010111,
    24'b111101111110011011011100,
    24'b111101011110010011011100,
    24'b111011001101110111010001,
    24'b001010110010010000100110,
    24'b000000000000000000000000,
    24'b000000000001100100111011,
    24'b000101110110000110111000,
    24'b000010110110011111001001,
    24'b000001000110001111010001,
    24'b000000110110011111010000,
    24'b000000110110010111010000,
    24'b000000100110010111010011,
    24'b000000000110011011010101,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000000110011111010010,
    24'b000000000110100011001101,
    24'b000001000110010011010001,
    24'b000001010110010011010010,
    24'b000101100101101110100011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b011000010101001101001011,
    24'b111100001110010011011011,
    24'b111011111110000111011001,
    24'b111100111110000111010101,
    24'b111100001110000011010011,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111011111110000111010110,
    24'b111011011101111111010100,
    24'b111100011110001011010111,
    24'b111100011110000011001110,
    24'b111000111101011011011010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000010000011010001101010,
    24'b000010010101111110111111,
    24'b000001100110100111010111,
    24'b000000010110011011001111,
    24'b000000110110010111010000,
    24'b000000110110010111010100,
    24'b000000000110011111010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010100,
    24'b000000010110010111010100,
    24'b000001010110010011010010,
    24'b000101000110001111000000,
    24'b000001110010101001011110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111100011110011011100000,
    24'b111010101110000011010111,
    24'b111100001110010011011001,
    24'b111100101110001011010100,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111011011101111011010000,
    24'b111011101110000011011011,
    24'b100011101000001110000010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000110000101101110101001,
    24'b000001010110100011001101,
    24'b000000000110011111010010,
    24'b000000010110100011010001,
    24'b000000110110011011001100,
    24'b000000010110011111001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100011001110,
    24'b000000110110011011001011,
    24'b000001010110001111010101,
    24'b000000110110010011001101,
    24'b000110010101011010010101,
    24'b000000000000110100101011,
    24'b000000000000000000000000,
    24'b110001111011111010111100,
    24'b111001111101110011010110,
    24'b111100001110001011011010,
    24'b111011111101111111010101,
    24'b111100111110000111011000,
    24'b111100101110000111011001,
    24'b111100101110000111011001,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000011011000,
    24'b111100111110000011011001,
    24'b111100111110000011011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100001110001011010111,
    24'b111101011110000111011000,
    24'b111010001110001111011001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000110010010101000110,
    24'b000101100110011110111011,
    24'b000001010110010111010101,
    24'b000000000110100011010010,
    24'b000000000110100011000111,
    24'b000000010110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001100,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111001101,
    24'b000000100110011111010010,
    24'b000000000110011111010011,
    24'b000001000110100011001010,
    24'b000000110110000111010000,
    24'b000011110110010111000010,
    24'b000001100010001001001001,
    24'b000000000000000000000000,
    24'b001110100011010000110010,
    24'b111100001110010111100000,
    24'b111100011110001011011011,
    24'b111100001110001011010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010110,
    24'b111100011110000011010110,
    24'b111100111110000111011010,
    24'b111011011110001111011010,
    24'b110001011011100110110111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001000010110001010100010,
    24'b000001100110000111001110,
    24'b000001100110011011001111,
    24'b000000000110101011010100,
    24'b000000000110011111010011,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001100,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001100,
    24'b000000100110011011010010,
    24'b000000100110010111010011,
    24'b000000100110101011000111,
    24'b000011110110110111010010,
    24'b000111110101101110100110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110011011100010010111110,
    24'b111100111110010111011101,
    24'b111100111110001011011001,
    24'b111100001110001011010101,
    24'b111100001110001011010101,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110001111010110,
    24'b111100011110001111011011,
    24'b111011111101111111011000,
    24'b111100001110001011011011,
    24'b001100000010101000100110,
    24'b000000000000000000000000,
    24'b000000010010001101010010,
    24'b000101110110101011001010,
    24'b000010010110001111001100,
    24'b000000010110011111010100,
    24'b000000000110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000010110011011010010,
    24'b000001000110010011010010,
    24'b000000000110101111000101,
    24'b000010010110001111000001,
    24'b000010110010100101011101,
    24'b000000000000000000000000,
    24'b001011000010100000101000,
    24'b111011011110001011011000,
    24'b111100011110000011010100,
    24'b111100011101111111010011,
    24'b111100001110001011010101,
    24'b111011111110001111010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111011101110000111011001,
    24'b111011101101111111011000,
    24'b111100001110000011011000,
    24'b101110111011001010101110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001000100110000110101101,
    24'b000010100110011011010000,
    24'b000001010110010011001111,
    24'b000000000110011011001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000001000110010111010000,
    24'b000000000110101111001010,
    24'b000101100110100010111001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101001011010001010100011,
    24'b111011011110001111010111,
    24'b111100101110000111010100,
    24'b111101001110000111010011,
    24'b111100011110001011010101,
    24'b111100001110001011010110,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100001110001011011001,
    24'b111100101110000111011001,
    24'b111100111110001011011001,
    24'b111011111110001111011101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000111000100101010000100,
    24'b000010000110010011001100,
    24'b000001000110010111010000,
    24'b000000000110011111010001,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111001110,
    24'b000000000110011111010001,
    24'b000000000110011011010100,
    24'b000000010110011011010000,
    24'b000000110110011011001100,
    24'b000000110110100011001111,
    24'b000110000101011110010111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111010101110001011011110,
    24'b111100011110010011011011,
    24'b111100101110000111010111,
    24'b111100111101111111010101,
    24'b111100101110000111010101,
    24'b111100101110000111010111,
    24'b111100111110000011011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100011110000111011000,
    24'b111100101110000111010111,
    24'b111101001110001011010111,
    24'b111011001101111111010111,
    24'b011011110110100001100100,
    24'b000000000000000000000000,
    24'b000000000001010000111111,
    24'b000100100110010111000001,
    24'b000000110110011111010001,
    24'b000000000110011111010011,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111001100,
    24'b000000000110011111010001,
    24'b000000000110011011010110,
    24'b000000010110011011010000,
    24'b000000100110011111001000,
    24'b000011000110010011001111,
    24'b000000110010110101011010,
    24'b000000000000000000000000,
    24'b010001000100000101000001,
    24'b111101011110010011010111,
    24'b111100001110010011011101,
    24'b111100001110000111011001,
    24'b111101001110000011010111,
    24'b111100111110000111010111,
    24'b111100111110000011011000,
    24'b111101001110000011011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111011000,
    24'b111100111110000111010111,
    24'b111100111110000011010100,
    24'b111011101110000011011000,
    24'b110110101101000011001011,
    24'b000000000000000000000000,
    24'b000000000001000000101111,
    24'b000110010101111110101011,
    24'b000000110110011011001100,
    24'b000000100110011011001101,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011011010001,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011011010000,
    24'b000000010110011011001110,
    24'b000011000110010010111101,
    24'b000000010001000100101100,
    24'b000000000000000000000000,
    24'b100110101001011110010101,
    24'b111101011110010011011001,
    24'b111100011110010111011010,
    24'b111011101110000111010101,
    24'b111101011110001111011001,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111011011101110011010100,
    24'b111011101110001011011011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000111010101011010010011,
    24'b000001110110100011001010,
    24'b000000100110011111010110,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110011011010001,
    24'b000000010110011011010000,
    24'b000000010110011011001110,
    24'b000100010101111110110001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110110001101000111001011,
    24'b111100001101111011010001,
    24'b111100111110010111011010,
    24'b111100001110001011010111,
    24'b111100001101111111010101,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000011011000,
    24'b111100001101111111010111,
    24'b111011111110000111011010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000011100011110101110100,
    24'b000010010110011111000110,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000110110011011001101,
    24'b000111110101111110100110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111011001110000011011000,
    24'b111101101110001111010110,
    24'b111011111101111111010101,
    24'b111100001110001011010111,
    24'b111100111110001011011000,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111011101101110111010101,
    24'b111100111110000111011001,
    24'b100000110111010001101110,
    24'b000000000000000000000000,
    24'b000000000001111001001100,
    24'b000010110110010010111111,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000010110011011001111,
    24'b000000100110011111010001,
    24'b000001010110010111001011,
    24'b001000100101001010001111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111100101110000111010111,
    24'b111101001110001011011000,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100011110001011010111,
    24'b111100011110001011010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100111110001011011010,
    24'b111100001101110111010011,
    24'b110100101100010010111110,
    24'b000000000000000000000000,
    24'b000000000000111100110011,
    24'b000011100110000110111100,
    24'b000000000110011111001110,
    24'b000000000110011111010001,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011011001111,
    24'b000000010110011011010010,
    24'b000001110110011011001101,
    24'b000110010011111101110011,
    24'b000000000000000000000000,
    24'b001010000010001000100001,
    24'b111100101110000011010101,
    24'b111100111110001011011011,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100001101111111010111,
    24'b111101011110001011011000,
    24'b110111111101010111001111,
    24'b000000000000000000000000,
    24'b000000000000101100101001,
    24'b000100100110001010111011,
    24'b000000000110011111001110,
    24'b000000000110011011010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111001111,
    24'b000000010110011111001111,
    24'b000000010110011011001111,
    24'b000010000110011111001100,
    24'b000011110011001001100101,
    24'b000000000000000000000000,
    24'b010100100100111001001100,
    24'b111100111110001111010110,
    24'b111011111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000011011000,
    24'b111100101110000111011001,
    24'b111100101110000111010110,
    24'b111000111101101011010010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000101010110001010111000,
    24'b000000100110011011010000,
    24'b000000010110011011010001,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010000,
    24'b000001010110011111010010,
    24'b000010010110011111001100,
    24'b000001100010110001011111,
    24'b000000000000000000000000,
    24'b011001100110001001011110,
    24'b111100101110001111010111,
    24'b111100101110001011010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011011000,
    24'b111001111101111111010110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000101000110001010110000,
    24'b000000100110010111010001,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010000,
    24'b000001010110011111010100,
    24'b000010010110011111001101,
    24'b000001100010100101011100,
    24'b000000000000000000000000,
    24'b011010000110001101100000,
    24'b111101001110001011011000,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111011111110001111010111,
    24'b111001101110000011010110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000101110110000110110000,
    24'b000000000110011011001111,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000100110100011010010,
    24'b000001000110011011010011,
    24'b000010010110011111001101,
    24'b000001110010110101011111,
    24'b000000000000000000000000,
    24'b010110110101010001010010,
    24'b111101001110000111011000,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100011110000011010110,
    24'b111100001110001011010111,
    24'b111100001110001111011000,
    24'b111001011101111111010100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000101000110000010110001,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000001010110011011010100,
    24'b000010000110011111001110,
    24'b000100010011101101101111,
    24'b000000000000000000000000,
    24'b001110010011001000110000,
    24'b111100101110000011010111,
    24'b111100011110000011010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111000011101101011010010,
    24'b000000000000000000000000,
    24'b000000000000100000101110,
    24'b000100100110000110110111,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000010110011111010000,
    24'b000001010110100011010001,
    24'b000001100110100011001101,
    24'b000111110101000010000101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111101001110000111010110,
    24'b111100101110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110001011011000,
    24'b111011111110000111010110,
    24'b111100001110000111010111,
    24'b110110111101010011001110,
    24'b000000000000000000000000,
    24'b000000000000110100110101,
    24'b000100000110010010111010,
    24'b000000000110011111010011,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111010010,
    24'b000000000110011111001111,
    24'b000000010110011111001100,
    24'b000000010110010011001001,
    24'b000111010101100110011011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111011111110001111011000,
    24'b111100101110001011010011,
    24'b111100001110001011010111,
    24'b111100001110001011011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100101110000111011000,
    24'b111011101110000011010111,
    24'b101010011010000010100000,
    24'b000000000000000000000000,
    24'b000000000001001101000100,
    24'b000010010110001011000100,
    24'b000000000110011111001011,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011111010001,
    24'b000000000110011111001111,
    24'b000000100110011111001101,
    24'b000000010110010111001100,
    24'b000111010101111010101011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111011001101111111011000,
    24'b111100011110000111010111,
    24'b111100001110001011011001,
    24'b111100001110001011011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100001101111111010111,
    24'b111011111110000011011001,
    24'b001111110011010100110101,
    24'b000000000000000000000000,
    24'b000011010010111101100010,
    24'b000010010110001111000111,
    24'b000000000110011111001100,
    24'b000000010110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000100110011111001110,
    24'b000000110110011011001111,
    24'b000101100101111110110101,
    24'b000000000000111000101110,
    24'b000000000000000000000000,
    24'b101111011011001010101000,
    24'b111011111110000011011010,
    24'b111100001110000111011001,
    24'b111100001110001011011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100111110001011011010,
    24'b111011101110000111011001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000111110100111010001000,
    24'b000010010110010011001001,
    24'b000000010110011011010010,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100011001110,
    24'b000000000110011111001110,
    24'b000000100110011111001111,
    24'b000000100110010011001111,
    24'b000100000110001110111110,
    24'b000000100001111001001000,
    24'b000000000000000000000000,
    24'b011100110110100101100001,
    24'b111011111110001011011010,
    24'b111100101110010011011011,
    24'b111011111110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000011010111,
    24'b111011111101111011010110,
    24'b111001011101011111010010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000110110101101110100011,
    24'b000001100110011111001100,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110100011001100,
    24'b000000000110011111001101,
    24'b000000010110011011010000,
    24'b000001010110100011010010,
    24'b000001110110011011000110,
    24'b000101010100101110000111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111011101110011011011101,
    24'b111011111110000111011000,
    24'b111100001110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000011011000,
    24'b111100111110001011011010,
    24'b101101111010110010100110,
    24'b000000000000000000000000,
    24'b000000000000110000111000,
    24'b000110000110010011000000,
    24'b000001000110100011010000,
    24'b000000010110011011001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110100011001100,
    24'b000000000110011011001101,
    24'b000000000110010111001111,
    24'b000001100110100111010011,
    24'b000000010110011011001110,
    24'b001000010110001010101110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110011111100100011000010,
    24'b111011111110001011011001,
    24'b111100101110001111011010,
    24'b111100011110000011010110,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110001011011001,
    24'b111100101110000111011000,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011011010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000011110010100101100010,
    24'b000011100110001111001010,
    24'b000000010110101011010101,
    24'b000000000110100011001101,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000001100110100111010000,
    24'b000000010110011111010101,
    24'b000101010110011011001001,
    24'b000001000001111001001011,
    24'b000000000000000000000000,
    24'b011000010101100001010111,
    24'b111010111101111011010101,
    24'b111100011110001111011001,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111011000,
    24'b111100111110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111011101110001111010110,
    24'b111100101110000011011001,
    24'b111101011110000011011000,
    24'b111100001110001011010110,
    24'b110111011101001011001100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000110100101001010011111,
    24'b000010000110001111001110,
    24'b000000010110011111010110,
    24'b000000110110011111010001,
    24'b000000010110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000100110011111010001,
    24'b000000010110100011010011,
    24'b000000010110011011010100,
    24'b000010110110010011001000,
    24'b000101010100101010001010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111011111110001111011101,
    24'b111100001110000111011000,
    24'b111100111110001111010110,
    24'b111100111110000111010101,
    24'b111100101110000111010110,
    24'b111100001110001011010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010011,
    24'b111100111110001011010001,
    24'b111100011110000111010110,
    24'b111011101110010011100000,
    24'b011011000110100001100100,
    24'b000000000000000000000000,
    24'b000000000001011100111110,
    24'b000110000110101011000001,
    24'b000001000110001011000111,
    24'b000000000110011111010011,
    24'b000000010110011011010001,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000100110011111010001,
    24'b000000100110100011010010,
    24'b000000000110011011010011,
    24'b000001010110010111010000,
    24'b000001110110001111001000,
    24'b000110000110001110110101,
    24'b000000100001001100110100,
    24'b000000000000000000000000,
    24'b011110010110111001101001,
    24'b111011111110001011011010,
    24'b111100011110000011010110,
    24'b111100101110001011010011,
    24'b111100011110001011010101,
    24'b111100001110001011010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111101001101111111011001,
    24'b111100011110000111010010,
    24'b111011111110000111010111,
    24'b111010001101101111011100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000100000100100110001100,
    24'b000000000110100111001011,
    24'b000000110110010111000101,
    24'b000000010110100011010000,
    24'b000000010110011011010001,
    24'b000000010110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010011,
    24'b000001110110011011010000,
    24'b000001110110010111001010,
    24'b000011000110010011000101,
    24'b000011000011110001110110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111011001110001111011110,
    24'b111011001101111111010011,
    24'b111100001110001011010110,
    24'b111100011110000011010101,
    24'b111100111110001011011010,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101101111111011001,
    24'b111100011110010011011011,
    24'b111011101110000011011000,
    24'b011010000101011101010111,
    24'b000000000000000000000000,
    24'b000000010001000000101110,
    24'b000110010110010110111011,
    24'b000000000110110011011000,
    24'b000000110110011011001001,
    24'b000000000110100011001101,
    24'b000000000110011011010001,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000100110011011010011,
    24'b000000100110011011010110,
    24'b000000010110011011001110,
    24'b000001110110011011001111,
    24'b000110100110010010111100,
    24'b000000000001010100111100,
    24'b000000000000000000000000,
    24'b010001110100000100111110,
    24'b111010111110000111011000,
    24'b111100001110001011010101,
    24'b111100101110000011011000,
    24'b111100101101111111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111001111,
    24'b111011101110000011011010,
    24'b111000101101001111001110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000101100100100010001010,
    24'b000010110110001111000010,
    24'b000000110110010011010100,
    24'b000000010110011011010000,
    24'b000000010110011011001101,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110010111010111,
    24'b000000100110011111010110,
    24'b000000010110100111010011,
    24'b000011100110101111001000,
    24'b000101000100101110010100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101111111011010110110000,
    24'b111110001110011011011110,
    24'b111101011110001111011100,
    24'b111100001110001011010010,
    24'b111100111110000111010111,
    24'b111100011110000111011000,
    24'b111100111110001011011000,
    24'b111100111110000111010101,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110001011011000,
    24'b111011101101111111010011,
    24'b111100111110001011010110,
    24'b111100001101101111001000,
    24'b111011001110001111010100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000100001101001001010,
    24'b000101010110001110111101,
    24'b000001100110011011001100,
    24'b000000110110010111010010,
    24'b000000010110011011010001,
    24'b000000010110011011001111,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010001,
    24'b000000100110010111010100,
    24'b000000000110011111010010,
    24'b000001000110010111001000,
    24'b000110000110001011000001,
    24'b000010000010101001010110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111001011110000111011000,
    24'b111011001110010011010111,
    24'b111101011101111011010111,
    24'b111100111110000111010110,
    24'b111100001110001011011001,
    24'b111100011110000011010110,
    24'b111101001110000011010101,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110001011010101,
    24'b111011011101110111010000,
    24'b111011011101110111011000,
    24'b011010100110010101011111,
    24'b000000000000000000000000,
    24'b000000000000101000101000,
    24'b000110000101011010100000,
    24'b000001110110011111001011,
    24'b000001100110101111010101,
    24'b000000000110010111001111,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011011001110,
    24'b000001000110010011010010,
    24'b000000000110001111001111,
    24'b000000110110100011010001,
    24'b000011010110011011001101,
    24'b000101110101110110110011,
    24'b000000000001001000110011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111001001101111111010101,
    24'b111110011101110011011000,
    24'b111100011110000111011000,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100111110001011011010,
    24'b111100111110001011011000,
    24'b111100111110000111010111,
    24'b111100101110000111011000,
    24'b111101001110010011011011,
    24'b101100011010011110100101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000101100100000101111101,
    24'b000010100110011111001000,
    24'b000000000110011011010000,
    24'b000000100110011111010001,
    24'b000000100110011111010001,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000010110011011010011,
    24'b000000100110010111010100,
    24'b000000100110011011010011,
    24'b000000000110010111001101,
    24'b000001110110101011001110,
    24'b000010000110100011001001,
    24'b000101110101000010010101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010100010100011001000110,
    24'b111010111110001011011001,
    24'b111100101110010111011101,
    24'b111100111110000011010101,
    24'b111100101110000011010110,
    24'b111100001110000111011010,
    24'b111100011110000111010111,
    24'b111100101110000111010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001101111011010100,
    24'b111101001110001011011000,
    24'b111101001110001111011001,
    24'b111100011110001111011100,
    24'b110011101100001010111101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000001010010100101011100,
    24'b000101000110001010111001,
    24'b000000110110010111001100,
    24'b000000000110011111010100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010100,
    24'b000000000110011111010010,
    24'b000000000110011111010000,
    24'b000000010110011011001100,
    24'b000000110110011011001101,
    24'b000001000110100011000011,
    24'b000011110110010011001110,
    24'b000100110100001010001010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010101000101011101011001,
    24'b111010111101111111011001,
    24'b111101111110000011010101,
    24'b111110001110010011011011,
    24'b111011001110000111011101,
    24'b111011111110000111010110,
    24'b111100101110000111010100,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110001011011000,
    24'b111100111110001011011000,
    24'b111100011101111111010100,
    24'b111101011110001111010110,
    24'b111100011101111111010011,
    24'b111101001110010011011100,
    24'b110010001011111010111011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000100001110000111111,
    24'b000100100110001010110101,
    24'b000000110110011111001101,
    24'b000000110110011011001011,
    24'b000000010110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110101011001100,
    24'b000000000110100011001110,
    24'b000001010110010111010010,
    24'b000001100110001111010011,
    24'b000001010110001111010000,
    24'b000000100110100011010001,
    24'b000011000110001111000011,
    24'b000100010011110001110010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010011110100010101000001,
    24'b111100101101101111001111,
    24'b111101111110000111011010,
    24'b111011001110001011011111,
    24'b111100001110001011010111,
    24'b111100101110001011010100,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110000011010110,
    24'b111100001110000011010110,
    24'b111101001110001111010101,
    24'b111100011110000011010000,
    24'b111101111110011011011000,
    24'b101110101010110110100101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001011100111111,
    24'b000110010101110110101111,
    24'b000010000110010111001000,
    24'b000000100110101111010010,
    24'b000000000110100011010001,
    24'b000000000110010111001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110011111010101,
    24'b000000010110011111010101,
    24'b000000100110011111001110,
    24'b000001000110011011001011,
    24'b000001100110010111001111,
    24'b000011110110001111000100,
    24'b000100000011111101111100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001010000010001100100110,
    24'b111010001101111111011011,
    24'b111100011110000011010110,
    24'b111110001110010111010111,
    24'b111101001110000111010011,
    24'b111100101110000111010111,
    24'b111100001110001011011001,
    24'b111100001110001011010101,
    24'b111100101110001011010011,
    24'b111101011110000111011000,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110001011010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100111110000011011001,
    24'b111100101110000111010110,
    24'b111100101110001011010101,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111011000,
    24'b111100101110000111011001,
    24'b111011111110000111011000,
    24'b111100111110001011010010,
    24'b111100101110001011010110,
    24'b111011011101111111011100,
    24'b111100011110001011011101,
    24'b111100001101110011011000,
    24'b111011101110001111010100,
    24'b100011001000011110000001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001101100111110,
    24'b000010000110000010110100,
    24'b000001100110010011000001,
    24'b000000010110011011001011,
    24'b000000000110011011001110,
    24'b000000010110100011001110,
    24'b000000010110100011001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010000,
    24'b000000110110100011010100,
    24'b000000110110010111001101,
    24'b000000010110011011010000,
    24'b000001110110101111010100,
    24'b000100110110000110111011,
    24'b000101000100011110001010,
    24'b000000000000101000101000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101011101010100010101000,
    24'b111010011101111111011010,
    24'b111011111101110111010011,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000111010100,
    24'b111100101110001011010101,
    24'b111100101110000011010110,
    24'b111100001110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100101110000111010111,
    24'b111100111110000111010110,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000111011001,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000011011000,
    24'b111101111101111011011010,
    24'b111101111101111111010100,
    24'b111101001110000111010101,
    24'b111100111110000011011001,
    24'b111100001110000011010001,
    24'b111011101101101111010010,
    24'b010000110011110000110110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000110001111101000100,
    24'b000100100110001110110011,
    24'b000010010110011011000111,
    24'b000001110110100011001111,
    24'b000000000110010111010001,
    24'b000000000110100011010110,
    24'b000000000110011011010011,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110100011001111,
    24'b000000000110011111001100,
    24'b000000010110100011010101,
    24'b000000110110100011010001,
    24'b000000000110011011001101,
    24'b000000000110011111010001,
    24'b000001000110010111010001,
    24'b000011100110010111001001,
    24'b000101010101001010010111,
    24'b000000000001010100111000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010100000100011000111110,
    24'b111001011101011111010000,
    24'b111100001110000111011010,
    24'b111011111101111011010100,
    24'b111101011110010011011010,
    24'b111100101110000111011000,
    24'b111100111110010011010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111101001110000011010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011011001,
    24'b111100001110001011011001,
    24'b111100001110001011011001,
    24'b111100001110001011010111,
    24'b111100111110000111010111,
    24'b111100111110000011010111,
    24'b111010101110010111010101,
    24'b111011111110010011011010,
    24'b111100111110000011011101,
    24'b111100111110001011100011,
    24'b100111001001010110010101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000010010011010101101010,
    24'b000101110110010110110110,
    24'b000001000110101011010000,
    24'b000000100110011011010000,
    24'b000000010110011011010010,
    24'b000000000110011111010101,
    24'b000000010110101011011000,
    24'b000000000110010111010011,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000000110011111001101,
    24'b000000000110100011010010,
    24'b000000000110100011010000,
    24'b000000000110100011001011,
    24'b000000010110100011001010,
    24'b000000100110011011001101,
    24'b000000100110011011001110,
    24'b000001100110011011000110,
    24'b000110110110001010101101,
    24'b000010100010101101010100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b011011000110010001100100,
    24'b111000111101100011010001,
    24'b111011111110000011011100,
    24'b111011111110000011011100,
    24'b111011011110000111010101,
    24'b111101111110001111011010,
    24'b111101001110000011010111,
    24'b111101001110000011010111,
    24'b111101001110000011010111,
    24'b111100111101111111010110,
    24'b111100111110000011010111,
    24'b111100111110000111011000,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100101110001111011001,
    24'b111011111110001011011001,
    24'b111011111110000111011000,
    24'b111011111101111011010101,
    24'b111100101101111111011001,
    24'b111100101110000111011011,
    24'b111010011110010111011011,
    24'b101011001010101110011110,
    24'b001011110010011000011111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001010000111000,
    24'b000011010101000010010111,
    24'b000001110110011111000001,
    24'b000000000110010111001100,
    24'b000000110110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011011010000,
    24'b000000110110011011001101,
    24'b000000010110011111001100,
    24'b000000000110011111001110,
    24'b000000000110010111001110,
    24'b000010000110011011001010,
    24'b000101010110010010111011,
    24'b000110010100111110010010,
    24'b000000000001011001000100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010101110100101101001101,
    24'b110001011011100110111001,
    24'b111011001110010011011001,
    24'b111101011110011011011100,
    24'b111011101101111111010100,
    24'b111100011110001011010111,
    24'b111100011110001011010111,
    24'b111100011110000111010111,
    24'b111100011110000111010111,
    24'b111100001110001011011001,
    24'b111100101110000111011001,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010101,
    24'b111100111110000011010100,
    24'b111100101110000111010101,
    24'b111011111110001111011010,
    24'b111011001110001011011000,
    24'b111011001101111011011000,
    24'b111001011101001011010000,
    24'b100101101000000110000101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000001100011000101011110,
    24'b000111000110000110110010,
    24'b000010000110011011001011,
    24'b000000100110100111001010,
    24'b000000100110011111010000,
    24'b000000010110100011010001,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011011010011,
    24'b000000100110011011001110,
    24'b000000010110011011010010,
    24'b000000000110011011010100,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000100110010011001101,
    24'b000001010110011011010000,
    24'b000000100110010111010110,
    24'b000001010110010011001111,
    24'b000110100110001110111010,
    24'b000110000011111001111101,
    24'b000000010001001000110111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010110010101011101010000,
    24'b101011001010011110011111,
    24'b110110111101001111001010,
    24'b111001111101111111010101,
    24'b111011001110010111011011,
    24'b111011001110010011011011,
    24'b111100001110000111011010,
    24'b111100001110000111011011,
    24'b111100011110000111011011,
    24'b111100011110000111011001,
    24'b111100011110001011011000,
    24'b111100011110000111010101,
    24'b111001001101011011001100,
    24'b110011011100010010111011,
    24'b011111000111010001101110,
    24'b001100010010101100101010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000100000101100,
    24'b000001110010001101011011,
    24'b000110010101101110101000,
    24'b000000110110001111000001,
    24'b000010010110011111010001,
    24'b000010000110001111001001,
    24'b000001010110100011001010,
    24'b000000000110011011010010,
    24'b000000000110011111001110,
    24'b000000000110011011010001,
    24'b000000010110011011010000,
    24'b000000010110011011001110,
    24'b000000000110011111001111,
    24'b000000000110011011010001,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000000110011111001111,
    24'b000000000110011111001101,
    24'b000000010110011011010000,
    24'b000000100110011011010010,
    24'b000001000110010111001110,
    24'b000001010110011111001010,
    24'b000001110110010111000101,
    24'b000110110110100011000000,
    24'b000101110100101010001100,
    24'b000001010001111101001011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001101010011000100101101,
    24'b010000110011111100111110,
    24'b010001110100010001000011,
    24'b010001010100001101000011,
    24'b001110110011110000111010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001010100110110,
    24'b000010110011100001101111,
    24'b000110010101101010101010,
    24'b000100010110010111000101,
    24'b000001000110000111001000,
    24'b000000110110010011001011,
    24'b000001010110011011010000,
    24'b000001100110100011010110,
    24'b000000110110011111010110,
    24'b000000010110100011010001,
    24'b000000000110011111001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001101,
    24'b000000000110011111010000,
    24'b000000010110011011010010,
    24'b000001000110011011010011,
    24'b000001000110011111001111,
    24'b000000000110110011001110,
    24'b000000010110110011001111,
    24'b000010110110011111001110,
    24'b000101110110001011000001,
    24'b000111110101111010101011,
    24'b000011100100100010000010,
    24'b000010100010100001010011,
    24'b000000000000111100110100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000101100101011,
    24'b000000000001110001000111,
    24'b000010100011010101101110,
    24'b000110010101001010011001,
    24'b000100000110010111000010,
    24'b000011100110100011001001,
    24'b000010000110101011001110,
    24'b000000000110010011001001,
    24'b000000000110100011001100,
    24'b000000010110011011001110,
    24'b000000110110010111010000,
    24'b000000100110011011010011,
    24'b000000110110011111010110,
    24'b000000010110011111010010,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100011001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010011,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011111001110,
    24'b000000000110100111001011,
    24'b000000000110100111001100,
    24'b000000000110010111010001,
    24'b000001000110010011010101,
    24'b000001110110010111000110,
    24'b000011010110001010111100,
    24'b000100110101110110101011,
    24'b000101100101011010011001,
    24'b000100000100011110000010,
    24'b000100000011111101111010,
    24'b000011110011100101110111,
    24'b000011100011100001101111,
    24'b000011110011100101101101,
    24'b000100000011110001110011,
    24'b000101100100001110000001,
    24'b000101010101000010011011,
    24'b000101100101100110101010,
    24'b000100110101111010110100,
    24'b000011010110001010111010,
    24'b000010000110010111000011,
    24'b000001010110010111001101,
    24'b000000110110010111001111,
    24'b000000110110011011001101,
    24'b000000010110011111001011,
    24'b000000110110011011001011,
    24'b000000110110011011001010,
    24'b000000110110011011001101,
    24'b000000010110010111010000,
    24'b000000010110011011010001,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110010111010100,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011111001111,
    24'b000000010110011011001101,
    24'b000000110110011011001011,
    24'b000000100110011011001011,
    24'b000000010110011011001010,
    24'b000000010110011011001001,
    24'b000000100110011111001010,
    24'b000001000110100111001101,
    24'b000001100110100111001011,
    24'b000001110110100011000110,
    24'b000001110110011111000011,
    24'b000001100110011011000001,
    24'b000001110110011111000100,
    24'b000001010110011011000101,
    24'b000001000110010011001000,
    24'b000001000110011011001110,
    24'b000000110110011111010000,
    24'b000000010110100111001101,
    24'b000000000110100011001101,
    24'b000000000110011111010001,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010001,
    24'b000000000110011011010011,
    24'b000000000110011011010100,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011001111,
    24'b000000010110011111001111,
    24'b000000010110011111010000,
    24'b000000010110011011010001,
    24'b000000100110011011010010,
    24'b000000010110011011010011,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110100011001101,
    24'b000000010110011111001111,
    24'b000000010110011111010000,
    24'b000000000110010111010000,
    24'b000000100110011111010001,
    24'b000000110110011011010001,
    24'b000000110110011111001110,
    24'b000000110110100011001110,
    24'b000001010110011111001111,
    24'b000001010110011011010000,
    24'b000000110110010111001101,
    24'b000000100110011111001100,
    24'b000000110110011011001111,
    24'b000000110110011111010011,
    24'b000000010110100011010101,
    24'b000000000110100011001111,
    24'b000000010110011111001110,
    24'b000000100110010111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010010,
    24'b000000010110011011010011,
    24'b000000010110011111010010,
    24'b000000010110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011111010001,
    24'b000000000110011011010011,
    24'b000000000110011011010010,
    24'b000000010110011011010011,
    24'b000000100110011111010100,
    24'b000000100110011011010011,
    24'b000000110110010111010010,
    24'b000001000110010111010000,
    24'b000001010110010111010010,
    24'b000000100110010111010010,
    24'b000000010110011011010011,
    24'b000000010110010111010011,
    24'b000000000110010111010000,
    24'b000000000110011111001101,
    24'b000000000110011111001011,
    24'b000000010110011011001110,
    24'b000000010110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000000110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000010110011111010011,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000100110010111010000,
    24'b000000100110010111010000,
    24'b000000000110011011010010,
    24'b000000000110011111010100,
    24'b000000010110011011010010,
    24'b000000010110011011001111,
    24'b000000010110011111001100,
    24'b000000000110100011001011,
    24'b000000000110011111001111,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000000110011111001100,
    24'b000000000110011111001101,
    24'b000000010110100011001111,
    24'b000000100110100111010010,
    24'b000000000110100111010010,
    24'b000000000110100011010011,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000010110100111010100,
    24'b000000000110100111010110,
    24'b000000010110011111010011,
    24'b000000000110011111010000,
    24'b000000010110100011001111,
    24'b000000010110100011001111,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000
};

assign mem = memory;

logic [23:0] memory_yellow [0:4899] = '{
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100011001100,
    24'b000000000110100011001110,
    24'b000000000110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000010110011011010010,
    24'b000000010110011011010000,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011001111,
    24'b000000000110011011001111,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000010110011111010010,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000100110010111001111,
    24'b000000100110010111010000,
    24'b000000100110010111010000,
    24'b000000100110010111010000,
    24'b000000100110010111001111,
    24'b000000010110100011001111,
    24'b000000010110100011001111,
    24'b000000000110011111001100,
    24'b000000010110100011001101,
    24'b000000000110011111001100,
    24'b000000000110011111001100,
    24'b000000000110011111001100,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011001111,
    24'b000000010110100011001111,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110100011010011,
    24'b000000000110100011010011,
    24'b000000010110011111010011,
    24'b000000010110011111010011,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011011010000,
    24'b000000010110011011010010,
    24'b000000000110011111010001,
    24'b000000010110100011010001,
    24'b000000010110100011010000,
    24'b000000010110100011001111,
    24'b000000000110011111001110,
    24'b000000000110011111001101,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000100110100011001110,
    24'b000000010110011011001111,
    24'b000000100110011111010011,
    24'b000000100110011011010100,
    24'b000000100110011011010101,
    24'b000000000110100011010011,
    24'b000000000110100011010010,
    24'b000000000110100011010000,
    24'b000000000110100011010000,
    24'b000000100110100011001111,
    24'b000000100110100011001111,
    24'b000000010110011111010001,
    24'b000000000110011111001101,
    24'b000000000110011111001101,
    24'b000000010110100111010000,
    24'b000000100110100111010011,
    24'b000001010110100111010100,
    24'b000000110110011111010011,
    24'b000000110110011111010100,
    24'b000000010110011111010011,
    24'b000000100110011111010100,
    24'b000000100110011111010100,
    24'b000000100110011111010001,
    24'b000000100110011111010010,
    24'b000000100110011111010010,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001101,
    24'b000000000110011011001011,
    24'b000000000110010111001110,
    24'b000000010110011011010010,
    24'b000000010110010111010100,
    24'b000000000110010011010100,
    24'b000000010110100011001111,
    24'b000000010110011111001110,
    24'b000001000110011111001101,
    24'b000001000110011011001011,
    24'b000001100110010011001010,
    24'b000001100110010011001001,
    24'b000001110110010111001001,
    24'b000001010110010011000101,
    24'b000001100110011011000100,
    24'b000001100110011011000110,
    24'b000001110110011011001001,
    24'b000001010110010111001001,
    24'b000001000110011011001010,
    24'b000001000110011011001101,
    24'b000001000110011011001111,
    24'b000000110110010111010000,
    24'b000000110110010111010001,
    24'b000000100110011111010001,
    24'b000000100110011111010001,
    24'b000001000110011011010001,
    24'b000000100110011111010001,
    24'b000000000110010111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000100110011011010001,
    24'b000000010110011011001111,
    24'b000000000110010011001110,
    24'b000000010110011011001111,
    24'b000001010110101111010100,
    24'b000001000110100011010011,
    24'b000001000110010111001101,
    24'b000001010110011011001010,
    24'b000010000110010111000101,
    24'b000011010110001011000001,
    24'b000100110110001110111100,
    24'b000101110110000110111001,
    24'b000101010101110110110001,
    24'b000100110101101010101101,
    24'b000100110101101110101010,
    24'b000100110101101110101000,
    24'b000100110101101110101010,
    24'b000101110101111110110011,
    24'b000100010110010110110111,
    24'b000010100110001010111000,
    24'b000010010110001010111111,
    24'b000010000110010111000011,
    24'b000001000110010011000111,
    24'b000001010110010111001111,
    24'b000001000110011111001111,
    24'b000000100110100011001110,
    24'b000000110110100011010011,
    24'b000000110110010111010001,
    24'b000000010110100011001111,
    24'b000000000110100011010011,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010000,
    24'b000000010110011111010011,
    24'b000000010110011011001101,
    24'b000000000110011011001010,
    24'b000000100110010111001101,
    24'b000000110110101011010000,
    24'b000001000110001111001100,
    24'b000100000110100011001101,
    24'b000010010110001011000000,
    24'b000100100110011011000111,
    24'b000110010110001010110101,
    24'b001000000101100110011101,
    24'b000101000011111001110110,
    24'b000010010010011101010110,
    24'b000000000001011100111011,
    24'b000000000000110100101011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001001100110111,
    24'b000000010001110101001001,
    24'b000010110011000001100110,
    24'b000110110101001110010100,
    24'b000110000101111010100110,
    24'b000101010101111110110001,
    24'b000100000110001111000100,
    24'b000001010110011011001010,
    24'b000000110110100111001011,
    24'b000001110110100111001111,
    24'b000000010110011111001100,
    24'b000000010110010111010100,
    24'b000000000110011111010001,
    24'b000000000110100011001100,
    24'b000000100110011111001111,
    24'b000000100110011011010001,
    24'b000000010110011011001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000110110010111001111,
    24'b000000010110011011010000,
    24'b000000110110011011001110,
    24'b000000100110100011001101,
    24'b000000100110011111001111,
    24'b000001000110100111001011,
    24'b000011100110010011000100,
    24'b001000010101111010101110,
    24'b001000010100110010001010,
    24'b000001010010010101010000,
    24'b000000000001001000110011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110101111011100101001110,
    24'b110110001011110001001100,
    24'b110110011011101101001110,
    24'b110110101011110001001111,
    24'b110101101011101001001110,
    24'b110101111011101101011000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000100001000100111000,
    24'b000100000011100001110101,
    24'b000111110101101110101101,
    24'b000101110110100011001010,
    24'b000010000110011011000110,
    24'b000001100110010111001111,
    24'b000001000110010011001101,
    24'b000001010110011111001100,
    24'b000000010110011011001001,
    24'b000000100110010111001100,
    24'b000000110110010111010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110100011001110,
    24'b000001000110100011001111,
    24'b000000000110011111010110,
    24'b000000000110100011011010,
    24'b000011010110000111000110,
    24'b000111100101110010110000,
    24'b000011110011101101111000,
    24'b000000000001010000111101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001010010000101100000101,
    24'b101111001010000000101101,
    24'b111100011100100100110111,
    24'b111110101100010100101111,
    24'b111111011100101100001101,
    24'b111111011100101000001010,
    24'b111111111100101000001100,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001100,
    24'b111111111100100100001100,
    24'b111111101100100100010001,
    24'b111111111100100100001111,
    24'b111111101100101100001010,
    24'b111110011100011100100111,
    24'b111100101100100100111000,
    24'b101111111010000100110001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000110000101111,
    24'b000001010010001101010100,
    24'b000110000100111010010110,
    24'b000100010110001110110111,
    24'b000001110110100011001001,
    24'b000000100110011111001010,
    24'b000000010110001011001101,
    24'b000000010110100011010101,
    24'b000001000110101111011000,
    24'b000000100110010011010010,
    24'b000000010110011011010000,
    24'b000000100110011111010001,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010000,
    24'b000000000110011111010000,
    24'b000000000110100011001100,
    24'b000010010110100011001000,
    24'b000011010110011011001001,
    24'b000100110101111010111001,
    24'b000100010011111001111100,
    24'b000000100001000100110101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100111111000001100110100,
    24'b111101001100101100011010,
    24'b111111011100101100001111,
    24'b111111111100100000001100,
    24'b111111111100100000010000,
    24'b111111111100100100001010,
    24'b111111011100101000001101,
    24'b111111111100100100001110,
    24'b111111111100100000001111,
    24'b111111111100100100010000,
    24'b111111111100100100010000,
    24'b111111111100100100001101,
    24'b111111111100101000001010,
    24'b111111111100100100001100,
    24'b111111001100101100001101,
    24'b111111111100100000010010,
    24'b111111111100011100010010,
    24'b111111001100011100001011,
    24'b111110111100101000001100,
    24'b111110111100100100010011,
    24'b111101101100011100101101,
    24'b100111011000000100111000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000001010010011001010111,
    24'b000101000101011110011111,
    24'b000011010110100011000001,
    24'b000001100110110111010011,
    24'b000001000110010011010001,
    24'b000010000110001011001011,
    24'b000001110110010111001000,
    24'b000000110110011011001110,
    24'b000000110110010111010000,
    24'b000000010110011011010000,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000010110100011010001,
    24'b000000010110011111010001,
    24'b000001010110010111001110,
    24'b000100100110010111000010,
    24'b000101110100111110010010,
    24'b000000000001010000111000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110001101010011000111100,
    24'b111111011100100000011001,
    24'b111111111100100000001010,
    24'b111111101100100100001111,
    24'b111111101100100000001101,
    24'b111111101100101000001110,
    24'b111111111100100100001110,
    24'b111111111100100100001010,
    24'b111111101100101100001101,
    24'b111111011100101100001011,
    24'b111111101100101000001011,
    24'b111111111100101000001101,
    24'b111111111100100100001110,
    24'b111111111100100100001101,
    24'b111111111100101000001100,
    24'b111111111100100100001110,
    24'b111111101100101000001100,
    24'b111111101100101000001100,
    24'b111111111100100100010000,
    24'b111111111100110000001110,
    24'b111111011100100000001110,
    24'b111111011100100100001110,
    24'b111111101100101000001110,
    24'b111111111100101000001101,
    24'b111111011100100000011101,
    24'b100001010110011100011100,
    24'b000000000000000000000000,
    24'b000000100000110000101001,
    24'b000010110011010001100111,
    24'b000110010110000110110011,
    24'b000011010110010111001011,
    24'b000001010110010011010000,
    24'b000000100110100011010010,
    24'b000000110110011011001110,
    24'b000000110110011011001110,
    24'b000000010110011011010000,
    24'b000000100110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011010000,
    24'b000000000110011011010011,
    24'b000000100110011111010011,
    24'b000000010110011011010000,
    24'b000000100110011111010010,
    24'b000000110110011111010101,
    24'b000001100110011111001010,
    24'b000010000110011111001101,
    24'b000110010110001010110100,
    24'b000011000011010101101011,
    24'b000000010000110000101001,
    24'b000000000000000000000000,
    24'b111000111100000001000010,
    24'b111111001100100000011010,
    24'b111111101100100100001111,
    24'b111111111100100100001110,
    24'b111111111100100100001110,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111101100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001110,
    24'b111111111100100100001100,
    24'b111111111100100100001101,
    24'b111111111100100100001100,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001110,
    24'b111111111100100100001100,
    24'b111111111100100100001101,
    24'b111111101100101000001100,
    24'b111111101100101000001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001100,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111110011100100000100000,
    24'b011110110110100000101001,
    24'b000000000000000000000000,
    24'b000000010001100000111110,
    24'b000110100101100110100010,
    24'b000011110110001011001001,
    24'b000010000110100111010000,
    24'b000000100110101111010011,
    24'b000000000110011011010010,
    24'b000000100110011011010001,
    24'b000001010110011111010010,
    24'b000000000110010111001101,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011010000,
    24'b000000000110011011010011,
    24'b000000000110011011010001,
    24'b000000000110100111001101,
    24'b000000010110011111001100,
    24'b000000100110010111010010,
    24'b000001010110010111000101,
    24'b000110100101101110101011,
    24'b000001010010001101010010,
    24'b000000000000000000000000,
    24'b010010110011010000010010,
    24'b111101101100100100100000,
    24'b111111001100101000001001,
    24'b111111111100100000001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111101100101000010000,
    24'b111100111100011100110110,
    24'b000000000000000000000000,
    24'b000000000000111100101011,
    24'b000101100100011101111101,
    24'b000101000110100110111111,
    24'b000001000110100011010000,
    24'b000001110110010011001101,
    24'b000010000110010111001011,
    24'b000000110110100111010001,
    24'b000000000110011011010000,
    24'b000000000110011111001101,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000100110011111010001,
    24'b000001000110010111001110,
    24'b000000000110011111010000,
    24'b000001010110010011010000,
    24'b000010010101110110111111,
    24'b000101000101011010011111,
    24'b000000110001011000111011,
    24'b000000000000000000000000,
    24'b011100000101011100011001,
    24'b111110101100101000010101,
    24'b111110001100011000010001,
    24'b111111111100101000001100,
    24'b111111011100101000001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111101100101100001101,
    24'b111111001100101100010001,
    24'b111101101100100000011011,
    24'b001010100001001000000101,
    24'b000000000000000000000000,
    24'b000011110011011101110101,
    24'b000100010110001111000001,
    24'b000010110110001111001010,
    24'b000000100110010011010000,
    24'b000000000110101011010100,
    24'b000000000110011111010010,
    24'b000000010110011011001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010011,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110010111001111,
    24'b000000010110010111010000,
    24'b000000100110011111010001,
    24'b000000100110011111010011,
    24'b000000100110011011010100,
    24'b000011000110010011001000,
    24'b000111000101111110011101,
    24'b000000000000110000110000,
    24'b000000000000000000000000,
    24'b111001011100000101000011,
    24'b111111001100100100001110,
    24'b111111111100011100010010,
    24'b111111111100100000001100,
    24'b111111011100101000001111,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111011100100100010000,
    24'b111111111100100100001011,
    24'b111111101100100100010001,
    24'b111111111100010100010110,
    24'b101011111001000000111011,
    24'b000000000000000000000000,
    24'b000011110011110001100111,
    24'b000100110110010010111101,
    24'b000000100110101011010010,
    24'b000000110110101011010101,
    24'b000000110110011011001100,
    24'b000000010110011111010000,
    24'b000000000110011111001110,
    24'b000000010110100011001111,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110010111010001,
    24'b000000110110100011010010,
    24'b000001000110011111001110,
    24'b000000100110011111001010,
    24'b000010000110010111000100,
    24'b000111010101111010101000,
    24'b000000100001001100111001,
    24'b000000000000000000000000,
    24'b111000001011101000111001,
    24'b111111011100101100001101,
    24'b111111001100011000001111,
    24'b111111111100100100010000,
    24'b111111001100101100000111,
    24'b111111111100101000001000,
    24'b111111011100101000001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001110,
    24'b111111111100101000001000,
    24'b111111111100100000001111,
    24'b111111011100100100001011,
    24'b111111011100101000010010,
    24'b101101101001010100111001,
    24'b000000000000000000000000,
    24'b000011010011111001101110,
    24'b000100010110011010111110,
    24'b000010010110010111001101,
    24'b000001010110010011010101,
    24'b000000010110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010011,
    24'b000000100110011011001111,
    24'b000001010110011111001111,
    24'b000010000110011011000111,
    24'b000110110110000010110010,
    24'b000000100001001100111001,
    24'b000000000000000000000000,
    24'b110111101011101000110111,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111101100101100001100,
    24'b111111011100101000010000,
    24'b111111111100100100001011,
    24'b111111101100100100010100,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111001100101100001101,
    24'b111111111100011100010000,
    24'b111111111100100000001110,
    24'b111110111100101100001100,
    24'b111111011100101100010000,
    24'b111111111100101000010010,
    24'b101000011000110000101111,
    24'b000000000000000000000000,
    24'b000110000100111110000011,
    24'b000100000110000011000100,
    24'b000001000110010011010010,
    24'b000000000110011111001111,
    24'b000000010110011111010101,
    24'b000000000110011011010010,
    24'b000000000110011111010001,
    24'b000000000110011111001110,
    24'b000000000110011111001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010010,
    24'b000000010110011011001111,
    24'b000000110110011011001101,
    24'b000000000110100011010100,
    24'b000001110110100111010000,
    24'b000001100110010011001000,
    24'b000101000110010010111101,
    24'b000001110010101101011101,
    24'b000000000000000000000000,
    24'b110111011011100001001110,
    24'b111111011100100000001011,
    24'b111111011100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111110011100100000010010,
    24'b010001000010111100010000,
    24'b000000000000000000000000,
    24'b000111000101101010100011,
    24'b000011110110011111001001,
    24'b000001100110011111010010,
    24'b000001100110011111010101,
    24'b000000010110010111010101,
    24'b000000010110011011010011,
    24'b000000010110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001100,
    24'b000000000110100011001011,
    24'b000000010110011111010000,
    24'b000000000110001111001011,
    24'b000011000110001010111000,
    24'b000100010100000001111101,
    24'b000000000000000000000000,
    24'b011010110101001000100000,
    24'b111111011100101000010101,
    24'b111111101100100000001101,
    24'b111111011100100100001111,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111001100100100001001,
    24'b111101111100100100011110,
    24'b000000000000000000000000,
    24'b000000100001100001000011,
    24'b000110110110000010110010,
    24'b000010010110100011001000,
    24'b000000100110001111010001,
    24'b000001000110011011010001,
    24'b000000110110010111010000,
    24'b000000100110010111010010,
    24'b000000010110011111010101,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010000,
    24'b000000010110011111010011,
    24'b000000010110011111010000,
    24'b000000110110011111010011,
    24'b000010010110010011001100,
    24'b000110010101101010100011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111111111100100000011101,
    24'b111111101100110000001110,
    24'b111111111100100000001010,
    24'b111111101100101000001010,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100101000010010,
    24'b111111101100101000001001,
    24'b111101011100010000111100,
    24'b000000000000000000000000,
    24'b000010000011010001100111,
    24'b000010110101111110111100,
    24'b000001100110100111010110,
    24'b000000000110011111010000,
    24'b000000110110011011001110,
    24'b000001000110010111001111,
    24'b000000010110011111010011,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110010111010100,
    24'b000000010110010111010101,
    24'b000001000110001111010001,
    24'b000101100110000110111100,
    24'b000001110010100101011111,
    24'b000000000000000000000000,
    24'b111011001100101001000010,
    24'b111111111100100000010010,
    24'b111111001100101100001111,
    24'b111111011100101000001110,
    24'b111111111100100000001111,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100101000001010,
    24'b111111101100100100001101,
    24'b111111101100101000001010,
    24'b100001100110101100100110,
    24'b000000000000000000000000,
    24'b000111000101101110100101,
    24'b000010010110011111001001,
    24'b000000000110011111010100,
    24'b000000010110011111010000,
    24'b000001000110011011001011,
    24'b000000010110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000110110011011001100,
    24'b000001010110001111010100,
    24'b000001100110001111001010,
    24'b000111000101011010010111,
    24'b000000010000111000101001,
    24'b010111010100010000100001,
    24'b111111011100101100001011,
    24'b111111111100100000001011,
    24'b111111011100101100001100,
    24'b111111101100100100010000,
    24'b111111111100100100001110,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001111,
    24'b111111101100100100001110,
    24'b111111011100101100001100,
    24'b111110011100100000100011,
    24'b000000000000000000000000,
    24'b000001010010010101001010,
    24'b000110010110011110111000,
    24'b000001010110010111010100,
    24'b000000010110100011010010,
    24'b000000110110011111001001,
    24'b000000000110011111010010,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000010110011111001111,
    24'b000000100110011111010011,
    24'b000000010110011011010011,
    24'b000000100110100011001001,
    24'b000000100110000111001010,
    24'b000100010110001011000010,
    24'b000001000010010101001000,
    24'b000000000000000000000000,
    24'b111101001100100000110011,
    24'b111111111100100100001110,
    24'b111111111100100000001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111101100101000001011,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001010,
    24'b111111111100011100010100,
    24'b111111101100101000001011,
    24'b111111101100101000001100,
    24'b101001011000010100101110,
    24'b000000000000000000000000,
    24'b001000010110000110100000,
    24'b000010010101110111001010,
    24'b000000110110011111001111,
    24'b000000110110100011010101,
    24'b000000000110100111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000010110011111001101,
    24'b000000100110011011010011,
    24'b000000110110010111010011,
    24'b000000010110100011000110,
    24'b000100110110110011010000,
    24'b000111100101101110100011,
    24'b000000000000000000000000,
    24'b010101100100001100011100,
    24'b111111001100100100010110,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111101100100000010001,
    24'b111111111100100100001010,
    24'b111111001100100000001101,
    24'b111101111100011100100101,
    24'b000000000000000000000000,
    24'b000000010010001101010110,
    24'b000110100110100011000110,
    24'b000010000110010111001001,
    24'b000000010110010111011000,
    24'b000000000110100011001100,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111001111,
    24'b000000010110011011010010,
    24'b000001000110010011010001,
    24'b000000010110100111000101,
    24'b000011100110000010111101,
    24'b000010100010101001011110,
    24'b000000000000000000000000,
    24'b111011111100100100111001,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111101100100100001111,
    24'b111111011100101000001100,
    24'b111111111100100100001101,
    24'b111111011100100100001101,
    24'b111111101100100000001011,
    24'b101110111001110100111100,
    24'b000000000000000000000000,
    24'b000111100110001110101000,
    24'b000011000110010111001100,
    24'b000000100110010111010001,
    24'b000000010110011011001110,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000001000110010111010000,
    24'b000000000110100111001100,
    24'b000110010110100010110100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111111101100100100010000,
    24'b111111111100100100001100,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001111,
    24'b111111011100101000001101,
    24'b111111111100100100001110,
    24'b111110111100110000001101,
    24'b111111111100100100001100,
    24'b111101101100100000101011,
    24'b000000000000000000000000,
    24'b000110100100011101111110,
    24'b000010110110001111001011,
    24'b000000110110011011001101,
    24'b000000000110011111010001,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110010111010100,
    24'b000000010110011011010001,
    24'b000000110110011011001100,
    24'b000001000110100011001100,
    24'b000111000101011010011010,
    24'b000000000000000000000000,
    24'b100111011000001000101101,
    24'b111111001100011000001101,
    24'b111111111100100100001110,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111101100100100010000,
    24'b111111001100101100001100,
    24'b111111101100100100010001,
    24'b111111001100100100010001,
    24'b000000000000000000000000,
    24'b000000000001010001000000,
    24'b000101010110010110111111,
    24'b000001000110011011010010,
    24'b000000010110100011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011011010001,
    24'b000000000110010111010101,
    24'b000000010110011011010000,
    24'b000000110110011111001000,
    24'b000011100110010111000111,
    24'b000001100010101101011110,
    24'b000000000000000000000000,
    24'b111110101100101100101111,
    24'b111111011100100100001000,
    24'b111111101100101000001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111001100101100001111,
    24'b111111111100100100001100,
    24'b111111111100100100010000,
    24'b111111111100011100001101,
    24'b111111111100100100001101,
    24'b111111011100101000001010,
    24'b110110011011101101010101,
    24'b000000010001001000101110,
    24'b000111100101110110101011,
    24'b000000100110100011001001,
    24'b000000100110010111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110011011010001,
    24'b000000010110011011010000,
    24'b000000010110011011001110,
    24'b000011100110001110111001,
    24'b000000010001001100110010,
    24'b000000000000000000000000,
    24'b111101101100110100011101,
    24'b111111011100011100001100,
    24'b111111111100100000001110,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100101000010000,
    24'b111101111100110000101001,
    24'b000000000000000000000000,
    24'b000111100101011010001101,
    24'b000010000110010111001100,
    24'b000000010110100011010010,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000110110011011001101,
    24'b000100110101111010101100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111111001100100000010001,
    24'b111111101100101000001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111001100101100010100,
    24'b000000000000000000000000,
    24'b000100000011101101110001,
    24'b000011110110011011000011,
    24'b000000010110011011010001,
    24'b000000010110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000001010110010111001010,
    24'b001000110101111110100010,
    24'b000000000000000000000000,
    24'b110000011001110100110011,
    24'b111111111100100100001001,
    24'b111111001100100100001011,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111011100101000010010,
    24'b000000000000000000000000,
    24'b000000000001111101001101,
    24'b000011110110001110111110,
    24'b000000100110011011001101,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110010111001111,
    24'b000000010110011011010000,
    24'b000001110110010011001010,
    24'b001001000101000110001010,
    24'b000000000000000000000000,
    24'b110000101001110100101111,
    24'b111111111100101000001011,
    24'b111111111100100100001110,
    24'b111111111100100100001110,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111001100100100001101,
    24'b001011010000111100000101,
    24'b000000000001001000110101,
    24'b000100010110000110110111,
    24'b000000010110100011001101,
    24'b000000000110011111010001,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011011001111,
    24'b000000000110010111010000,
    24'b000010000110011011001011,
    24'b000110100100000101110011,
    24'b000000000000000000000000,
    24'b111100011100100000110110,
    24'b111111111100101000001000,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100010000,
    24'b111110111100101000001101,
    24'b111011101100011100111110,
    24'b000000000000110000101110,
    24'b000101010110000110111001,
    24'b000000100110011011001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000010110011111001111,
    24'b000000010110011011001111,
    24'b000010000110011011001010,
    24'b000011100011000101100101,
    24'b000000000000000000000000,
    24'b111101011100100000101110,
    24'b111111111100100000001100,
    24'b111111011100101000001101,
    24'b111111111100100100001110,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111101100100100001111,
    24'b111111001100101000000011,
    24'b111101101100011100111001,
    24'b000000000000101000101100,
    24'b000101110110001010110010,
    24'b000000110110010111010000,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000010110011111001111,
    24'b000001010110100011010000,
    24'b000010110110011111001010,
    24'b000010000010101101011110,
    24'b000000000000000000000000,
    24'b111100101100100100101110,
    24'b111111111100100000001101,
    24'b111111101100101000001011,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111101100100100001101,
    24'b111111011100110100001011,
    24'b111101011100011000111100,
    24'b000000000000000000000000,
    24'b000101110110000110110010,
    24'b000000100110011011001110,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010000,
    24'b000001010110011111010010,
    24'b000011000110011011001011,
    24'b000001100010101101011010,
    24'b000000000000000000000000,
    24'b111100101100100100110000,
    24'b111111111100100000001111,
    24'b111111001100101100001100,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111101100100100001101,
    24'b111111101100101100001110,
    24'b111100111100010101000001,
    24'b000000000000000000000000,
    24'b000101110110000010101111,
    24'b000000010110011111001110,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000010110011111010010,
    24'b000001010110011111010011,
    24'b000011010110011011001011,
    24'b000010010010101101100011,
    24'b000000000000000000000000,
    24'b111100111100100100101101,
    24'b111111111100100100001101,
    24'b111111111100100100001111,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100011100001011,
    24'b111100001100100100110111,
    24'b000000010000011000101001,
    24'b000110000101111010110000,
    24'b000000010110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010001,
    24'b000001000110011011010010,
    24'b000010110110011011001011,
    24'b000100000011100101110011,
    24'b000000000000000000000000,
    24'b111100011100100100110100,
    24'b111111111100101000001010,
    24'b111111111100011100010000,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100011100001101,
    24'b111010001100011101000100,
    24'b000000000000101000110011,
    24'b000101110101111110110110,
    24'b000000100110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010011,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000010110011111001111,
    24'b000001010110100011010000,
    24'b000001110110011011001000,
    24'b000111000101000110000010,
    24'b000000000000000000000000,
    24'b110001001001110100101110,
    24'b111111001100101100001011,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111011100101000001100,
    24'b111111011100010100001111,
    24'b001011000001001000000101,
    24'b000000000001000000110100,
    24'b000101000110001010111001,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111001111,
    24'b000000010110011111001100,
    24'b000000100110010111000110,
    24'b000111110101100010011000,
    24'b000000000000000000000000,
    24'b110000111001110100110100,
    24'b111111001100101100001001,
    24'b111111011100100100001111,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111101100101000001110,
    24'b001010100001001100000110,
    24'b000000000001010101000011,
    24'b000011000110001010111110,
    24'b000000000110100011001100,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011111001111,
    24'b000000100110011111001101,
    24'b000000100110010111001010,
    24'b000111010101111010101011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111111101100100100010100,
    24'b111111101100101100001111,
    24'b111111111100100100001100,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001110,
    24'b111111101100100100010011,
    24'b000000000000000000000000,
    24'b000011100010111101100110,
    24'b000011000110001011000100,
    24'b000000000110011111001101,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000100110011111001111,
    24'b000000100110011111001100,
    24'b000101010110000010110101,
    24'b000000000001000000110001,
    24'b000000000000000000000000,
    24'b111111001100100100010101,
    24'b111111001100011100001011,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001100,
    24'b111110011100110000010000,
    24'b000000000000000000000000,
    24'b000111110100111010001011,
    24'b000011000110001011000110,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011001111,
    24'b000000000110011111001110,
    24'b000000100110011111001111,
    24'b000000100110010111001101,
    24'b000100000110001110111011,
    24'b000000100010000001000110,
    24'b000000000000000000000000,
    24'b111101011100110000011101,
    24'b111111111100100000010000,
    24'b111111111100100100001110,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100000001100,
    24'b110101111011001001001101,
    24'b000000000000000000000000,
    24'b000111100101101110011100,
    24'b000010100110010111001100,
    24'b000000010110010111010100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111001110,
    24'b000000010110100011001101,
    24'b000000000110011011001101,
    24'b000000010110010111001111,
    24'b000001000110100011010010,
    24'b000011010110011111000011,
    24'b000101010100110010000100,
    24'b000000000000000000000000,
    24'b101000001000010100110010,
    24'b111111001100011100001101,
    24'b111111111100100100001110,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111011100101100001101,
    24'b000000000000000000000000,
    24'b000000000000101000110111,
    24'b000110110110010010111011,
    24'b000001010110011111001110,
    24'b000000010110011011001100,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111001110,
    24'b000000000110011111001100,
    24'b000000000110011011001101,
    24'b000000000110010011001110,
    24'b000001010110101011010100,
    24'b000001010110011011001001,
    24'b000111010110001110110000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111110101100100100001111,
    24'b111111111100100000001110,
    24'b111111111100100100001100,
    24'b111111111100100100001110,
    24'b111111111100100100001100,
    24'b111111111100100100001100,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001110,
    24'b111101111100011100110000,
    24'b000000000000000000000000,
    24'b000011100010100001100001,
    24'b000100000110001011001000,
    24'b000000100110101111010010,
    24'b000000110110011011010001,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000001010110100111010010,
    24'b000000100110100011010001,
    24'b000101100110011011000110,
    24'b000001010001110001001010,
    24'b000000000000000000000000,
    24'b111100111100100000111001,
    24'b111111101100100100010000,
    24'b111111111100101000001011,
    24'b111111101100101000001110,
    24'b111111111100100100001101,
    24'b111111101100100100001111,
    24'b111111111100101000001010,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111101100101000001100,
    24'b111111111100100000001011,
    24'b111111011100100100010010,
    24'b111111111100101000001010,
    24'b111111001100100100010010,
    24'b110000011001110000111010,
    24'b000000000000000000000000,
    24'b000110110101000010011100,
    24'b000010000110001011001010,
    24'b000000110110010111010110,
    24'b000001010110011011010001,
    24'b000000010110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000100110011111010001,
    24'b000000110110011111010100,
    24'b000000010110011111001110,
    24'b000011100110001011001000,
    24'b000101110100101010001100,
    24'b000000000000000000000000,
    24'b010101100100010000011010,
    24'b111110111100101000010010,
    24'b111111101100101000001111,
    24'b111111111100100100010000,
    24'b111111001100101100001100,
    24'b111111101100100000010100,
    24'b111111111100100100001001,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111011100100100001111,
    24'b111111111100101000000111,
    24'b111111001100101000010011,
    24'b111111011100101000001010,
    24'b111110101100101000011100,
    24'b000000000000000000000000,
    24'b000000010001011101000001,
    24'b000110010110100010111111,
    24'b000000100110010011000110,
    24'b000000000110011111010010,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000100110011111010001,
    24'b000000100110100011010010,
    24'b000000110110010111010011,
    24'b000000010110011111001110,
    24'b000010010110001111001001,
    24'b000111010110001110110011,
    24'b000000110001001100110110,
    24'b000000000000000000000000,
    24'b111101011100011100110100,
    24'b111111011100101000001110,
    24'b111111111100100000001100,
    24'b111110111100101100001100,
    24'b111111101100100100001101,
    24'b111111111100100000001111,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001100,
    24'b111111111100100000010100,
    24'b111111011100101000001101,
    24'b111111111100011100001111,
    24'b101001011000000100110010,
    24'b000000000000000000000000,
    24'b000100110100100010001010,
    24'b000000100110010011000101,
    24'b000000100110011011000100,
    24'b000000000110100011010000,
    24'b000000000110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000110110010111010000,
    24'b000000110110100011010000,
    24'b000001010110010111001010,
    24'b000100000110001111000001,
    24'b000011100011110101110111,
    24'b000000000000000000000000,
    24'b010111000100011000100001,
    24'b111111111100101000001010,
    24'b111111011100101100001100,
    24'b111111111100100100001111,
    24'b111111111100011100001101,
    24'b111110111100110000001100,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100101000001011,
    24'b111111111100101000001000,
    24'b111110111100011100011011,
    24'b000000000000000000000000,
    24'b000000000001001100101111,
    24'b000111000110010010111000,
    24'b000001000110101111010010,
    24'b000000100110011111000111,
    24'b000000010110100011001101,
    24'b000000100110011011010010,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010001,
    24'b000001010110011011010111,
    24'b000000000110100011001011,
    24'b000001100110010111001111,
    24'b000110110110001110111101,
    24'b000000000001011100111110,
    24'b000000000000000000000000,
    24'b111011101100100101000011,
    24'b111110111100100000010001,
    24'b111111111100100100001101,
    24'b111111111100100100001010,
    24'b111111001100101100001111,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001111,
    24'b111111111100101000001100,
    24'b111111001100101000010010,
    24'b100011000111001000100100,
    24'b000000000000000000000000,
    24'b000101110100011110001000,
    24'b000011010110001111000000,
    24'b000000100110001111010101,
    24'b000000010110011011001111,
    24'b000000110110011011001101,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010011,
    24'b000000010110010111010110,
    24'b000000100110011111011000,
    24'b000001000110101011010011,
    24'b000100000110101011000101,
    24'b000101010100101110010000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111101111100101100011101,
    24'b111111101100100000001111,
    24'b111110111100100100001101,
    24'b111111101100100000001100,
    24'b111111111100100100001110,
    24'b111111111100101000001100,
    24'b111111111100100000001110,
    24'b111111111100100100001010,
    24'b111111111100100100001111,
    24'b111111111100101000001100,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100000010001,
    24'b111111111100100100001101,
    24'b111111001100101100001011,
    24'b111111111100100100001100,
    24'b111111111100100000001111,
    24'b111111111100011100001111,
    24'b111111001100011000001111,
    24'b111111111100101000001100,
    24'b111011101100011100111111,
    24'b000000000000000000000000,
    24'b000000110001101001000110,
    24'b000101100110001010111110,
    24'b000001100110010111001110,
    24'b000000100110010111010101,
    24'b000000010110011011010001,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010001,
    24'b000000100110010111010100,
    24'b000000000110011111010001,
    24'b000001100110010011000100,
    24'b000110110110001010111101,
    24'b000010000010100101011100,
    24'b000000000000000000000000,
    24'b011101000101101000100000,
    24'b111111101100100100011100,
    24'b111111111100100100001010,
    24'b111111101100101100001100,
    24'b111111011100101000001101,
    24'b111111011100101000001101,
    24'b111111111100100100010010,
    24'b111111111100100100001101,
    24'b111111111100100100001100,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111011100101000001101,
    24'b111111111100100100001100,
    24'b111111011100101000001101,
    24'b111111011100101100001011,
    24'b111111011100101000001101,
    24'b111111111100101000000110,
    24'b111111001100110000010110,
    24'b001011010001111000001110,
    24'b000000100000101000101010,
    24'b000110010101011010011111,
    24'b000010110110011111001100,
    24'b000001100110101111010101,
    24'b000000000110010111001111,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001101,
    24'b000000110110011011001100,
    24'b000001000110010011010010,
    24'b000000000110001011010001,
    24'b000001000110011111010001,
    24'b000011110110010011001101,
    24'b000110000101110110101101,
    24'b000000000001011000110100,
    24'b000000000000000000000000,
    24'b110110111011100101001110,
    24'b111111111100100000001010,
    24'b111111001100101000010010,
    24'b111111011100101100001101,
    24'b111111101100101000001101,
    24'b111111101100101000001110,
    24'b111111101100101000001100,
    24'b111111111100100100001110,
    24'b111111111100100100001100,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111001100101100001011,
    24'b111111111100100100001100,
    24'b111111111100100100001101,
    24'b111111101100101000001101,
    24'b111111011100101000001110,
    24'b111111011100101000001110,
    24'b111111111100100100010110,
    24'b100101010111110100111011,
    24'b000000000000000000000000,
    24'b000101100100000101111001,
    24'b000011000110011111000001,
    24'b000000000110011011010010,
    24'b000000100110011111010001,
    24'b000000100110011111010001,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000010110011011010011,
    24'b000001000110010011010101,
    24'b000000010110011011010100,
    24'b000000000110011011001111,
    24'b000010000110100111001110,
    24'b000011000110011011000100,
    24'b000110000101000110010111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111000111011100100110010,
    24'b111110111100101000001111,
    24'b111111111100100000010101,
    24'b111111111100100100001001,
    24'b111111101100011100010011,
    24'b111111011100101100001100,
    24'b111111111100100000010010,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001100,
    24'b111111011100101000001101,
    24'b111111011100101000001101,
    24'b111111111100011000010001,
    24'b111111011100101100001100,
    24'b111111111100100000010010,
    24'b101001101000101000110000,
    24'b000000000000000000000000,
    24'b000010000010100101011001,
    24'b000101000110001010110111,
    24'b000000110110010011001101,
    24'b000000100110011111010011,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110010111010101,
    24'b000000010110010111010100,
    24'b000000010110011111010001,
    24'b000000000110011011001100,
    24'b000001000110011011001011,
    24'b000001110110100011000010,
    24'b000100000110001111001001,
    24'b000100110100001010000101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110111111011101000110110,
    24'b111111001100110100001110,
    24'b111111111100100000001100,
    24'b111111111100100100001010,
    24'b111111011100101100001100,
    24'b111111011100101100001100,
    24'b111111111100100100001100,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100000010000,
    24'b111111011100101000001011,
    24'b111111101100100100001110,
    24'b111111011100101100001100,
    24'b111111001100101100010101,
    24'b101100111001010000111101,
    24'b000000000000000000000000,
    24'b000000100001111001000010,
    24'b000110000110000010110010,
    24'b000001100110011111000111,
    24'b000001000110011011001011,
    24'b000000110110010111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100011001110,
    24'b000000000110100111001101,
    24'b000000010110011011001110,
    24'b000000110110011011010001,
    24'b000001100110001111010010,
    24'b000000010110010011001111,
    24'b000001100110011111010010,
    24'b000100010110000110111111,
    24'b000100010011110101110001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111010001100000000111101,
    24'b111110101100101000001101,
    24'b111111011100011000001111,
    24'b111111011100100100010001,
    24'b111111011100101100001100,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100011100001110,
    24'b111111011100101000001101,
    24'b111111011100101000001110,
    24'b111111111100011100010010,
    24'b101100001001000000111001,
    24'b000000000000000000000000,
    24'b000000010001010100111101,
    24'b000110110101110110101010,
    24'b000001110110010011001000,
    24'b000000110110101111010010,
    24'b000000000110100111001111,
    24'b000000110110010111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011111010101,
    24'b000000010110011111010101,
    24'b000001000110011111001011,
    24'b000000110110010011001100,
    24'b000001100110010111001111,
    24'b000100110110001010111111,
    24'b000100100011111101111011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b011110110101011000011100,
    24'b111110101100100000010110,
    24'b111111111100100100001010,
    24'b111110111100011000001100,
    24'b111111111100100100001100,
    24'b111111111100100100001110,
    24'b111111011100100100010010,
    24'b111111101100101000001101,
    24'b111111111100100100001100,
    24'b111111011100101100001100,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111011100101000001110,
    24'b111111011100101000001101,
    24'b111111111100100000010001,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111011100100100010001,
    24'b111111111100100100001101,
    24'b111111111100100000001100,
    24'b111111101100101000001100,
    24'b111111001100101100001100,
    24'b111111111100100100001100,
    24'b111111101100011100001011,
    24'b111111101100101000001010,
    24'b111110011100100100011111,
    24'b001101000001011000000110,
    24'b000000000000000000000000,
    24'b000000100001110001000001,
    24'b000011100110000110110000,
    24'b000010010110001110111111,
    24'b000000110110010111001010,
    24'b000000000110011011001110,
    24'b000000010110100011001110,
    24'b000000000110011111001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000110110100011010100,
    24'b000000010110010111010001,
    24'b000000000110011011010011,
    24'b000010100110101011010001,
    24'b000101100110000010110110,
    24'b000101010100011010001001,
    24'b000000010000111000101011,
    24'b000000000000000000000000,
    24'b010011100011010100010001,
    24'b111101111100101000100100,
    24'b111111101100101000010001,
    24'b111111011100101100001010,
    24'b111111011100100100010001,
    24'b111111111100100000001101,
    24'b111111111100100000001100,
    24'b111111111100011100001110,
    24'b111111111100011100010001,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111101100100100001110,
    24'b111111111100101000001010,
    24'b111111111100100100001110,
    24'b111111111100101000001001,
    24'b111111111100100100001101,
    24'b111111111100101000001001,
    24'b111111101100101000001100,
    24'b111111111100100000010001,
    24'b111111111100100000001101,
    24'b111111111100100000001111,
    24'b111111101100100100010000,
    24'b111111011100011100010010,
    24'b111011111100100000111000,
    24'b001010100001101000001001,
    24'b000000000000000000000000,
    24'b000001010010000001001111,
    24'b000110000110010010110011,
    24'b000010110110010111000100,
    24'b000010010110100011001110,
    24'b000000010110010111010011,
    24'b000000000110011111010111,
    24'b000000000110011011010100,
    24'b000000010110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000010110100011001111,
    24'b000000000110011111001110,
    24'b000000010110011111010101,
    24'b000000110110100011010100,
    24'b000000000110011011001110,
    24'b000000010110100011010010,
    24'b000001010110010111001101,
    24'b000100000110001111001000,
    24'b000110100100111110011010,
    24'b000000000001100000110101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111001011011111101000001,
    24'b111111001100100100011000,
    24'b111111101100100100001101,
    24'b111111001100101100001110,
    24'b111111001100101100001101,
    24'b111111011100101100001011,
    24'b111111101100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100000010010,
    24'b111111111100100100001011,
    24'b111111011100100000010111,
    24'b111111011100101100001100,
    24'b111111111100100100001101,
    24'b111111111100100000001101,
    24'b111111111100100000010010,
    24'b111110111100101100001101,
    24'b111111101100101000001000,
    24'b111111111100100100001111,
    24'b111101111100101000100000,
    24'b100001100110010100100110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000010110011001101101101,
    24'b000110010110010110110101,
    24'b000010000110100111001101,
    24'b000001000110011011001110,
    24'b000000010110010111010001,
    24'b000000000110011111010101,
    24'b000000010110101011011001,
    24'b000000000110010111010011,
    24'b000000000110010111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000010110100011010010,
    24'b000000010110011111001110,
    24'b000000010110100011001011,
    24'b000000010110100011001011,
    24'b000000110110011011001101,
    24'b000001000110011011001111,
    24'b000001100110011011000110,
    24'b001000010110000110101101,
    24'b000010110010100101010110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110011001010100000111000,
    24'b111111001100100100011000,
    24'b111111101100100000001111,
    24'b111111001100100100001010,
    24'b111111111100011100010011,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001110,
    24'b111111111100101000001010,
    24'b111111101100101100001011,
    24'b111111101100101100001110,
    24'b111111011100100000010000,
    24'b111111001100101000001001,
    24'b111111011100101100001110,
    24'b111111101100100000001001,
    24'b111110011100100100011100,
    24'b100010100110110000011011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001011000111110,
    24'b000011110100111110010101,
    24'b000011010110010011000011,
    24'b000000110110010111000111,
    24'b000000000110100111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000010110011011001111,
    24'b000000110110011011001101,
    24'b000000010110011011001101,
    24'b000000000110011111001100,
    24'b000000010110010111001011,
    24'b000010110110010111001000,
    24'b000101000110001110111100,
    24'b000101010100111010001101,
    24'b000000000001011101000100,
    24'b000000000000101000101100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110000101001111000110001,
    24'b111110101100101000011100,
    24'b111111011100101100010000,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100100001110,
    24'b111111111100100100001110,
    24'b111111111100100100001101,
    24'b111111101100011100010001,
    24'b111110011100110000000110,
    24'b111110011100101100011000,
    24'b111110101100101100011100,
    24'b101000101000001100110001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000100100101000,
    24'b000001100011000001100000,
    24'b001000000110000110101100,
    24'b000011010110010011001011,
    24'b000000000110110011001011,
    24'b000000010110100011001100,
    24'b000000010110100011001110,
    24'b000000000110011011010011,
    24'b000000000110011111001111,
    24'b000000000110011111001100,
    24'b000000000110011111001101,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011011010011,
    24'b000000000110011111001110,
    24'b000000000110011011010010,
    24'b000000000110011011010100,
    24'b000000010110010111010011,
    24'b000000000110011111010001,
    24'b000000010110100011010000,
    24'b000000010110001111010001,
    24'b000000110110011111001110,
    24'b000000110110010111010011,
    24'b000010110110001111001100,
    24'b000111000110001010110110,
    24'b000101010100000101111011,
    24'b000000010001001000111100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001011110001110000000101,
    24'b110000101010001000101101,
    24'b111100111100100000110101,
    24'b111110111100100000011101,
    24'b111111111100101000001100,
    24'b111111111100100100010000,
    24'b111111111100100100001110,
    24'b111111101100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100000001100,
    24'b111111111100100100001101,
    24'b111111111100100100001101,
    24'b111111111100100000010001,
    24'b111111101100100100001100,
    24'b111110011100011100100011,
    24'b111100111100101000111000,
    24'b101111111010001000110001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000101000110000,
    24'b000001100010010101011110,
    24'b000101110101100110100011,
    24'b000010000110000110111101,
    24'b000010010110100011010000,
    24'b000001000110011011001011,
    24'b000001110110011111001001,
    24'b000000110110010111010001,
    24'b000000100110010011010010,
    24'b000000000110011011010100,
    24'b000000010110011011010000,
    24'b000000010110011011001110,
    24'b000000000110011111001111,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000100110100111010010,
    24'b000000000110011111010000,
    24'b000000010110011011001101,
    24'b000000010110011011010010,
    24'b000000100110011011010010,
    24'b000001000110010111001110,
    24'b000010000110011011001000,
    24'b000010110110001111000001,
    24'b000111110110011110111010,
    24'b000110010100101110001011,
    24'b000001010010000001001011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001100100001011100000000,
    24'b110110011011110001001101,
    24'b110111001011101001001110,
    24'b110111001011101001001110,
    24'b110110101011100001001101,
    24'b110110101011100001001100,
    24'b110110101011100101001101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001011000111001,
    24'b000011010011100001101111,
    24'b000111000101100110100101,
    24'b000101000110010011000001,
    24'b000001000110000011000011,
    24'b000000100110001111001010,
    24'b000001000110100011001111,
    24'b000001100110100011010100,
    24'b000000110110011111010110,
    24'b000000010110011111010010,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011011001101,
    24'b000000000110011011010010,
    24'b000000000110011011010100,
    24'b000000010110011011010010,
    24'b000000110110011011001110,
    24'b000000010110110111010000,
    24'b000000110110110011001111,
    24'b000011100110011111001001,
    24'b000110010110000110111010,
    24'b001000100101111010101001,
    24'b000011100100010110000100,
    24'b000001100010100101011010,
    24'b000000000001000000110010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000100100101110,
    24'b000001000010001101001110,
    24'b000011100011100001110001,
    24'b000110110100111010011110,
    24'b000101100110001110111101,
    24'b000100100110011111000101,
    24'b000010100110100011001010,
    24'b000000000110001111001001,
    24'b000000000110011111001110,
    24'b000000010110011111001101,
    24'b000000110110011011001110,
    24'b000000110110011011010010,
    24'b000000110110100011010100,
    24'b000000010110011111010010,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010011,
    24'b000000000110011011010100,
    24'b000000000110011011010011,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000010110100111001110,
    24'b000000100110100011001101,
    24'b000001000110010111001101,
    24'b000001100110010011010000,
    24'b000010100110001111000100,
    24'b000100000110001010110110,
    24'b000101000101111010100101,
    24'b000101110101011010010110,
    24'b000100100100011010000110,
    24'b000100100011111101110110,
    24'b000100010011100101110101,
    24'b000011110011011101101111,
    24'b000100010011100101101111,
    24'b000100000011101101110010,
    24'b000101100100001001111111,
    24'b000110000101000010011000,
    24'b000110010101100110101001,
    24'b000101010101111110101100,
    24'b000011010110001110111001,
    24'b000010000110011110111100,
    24'b000001010110011011001001,
    24'b000001000110010111001111,
    24'b000000100110010111001101,
    24'b000000010110011011001101,
    24'b000000110110011011001100,
    24'b000000100110011011001100,
    24'b000000110110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011010001,
    24'b000000010110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010100,
    24'b000000100110010111010001,
    24'b000000100110010111010000,
    24'b000000010110011011010001,
    24'b000000010110011111010001,
    24'b000000000110011111001110,
    24'b000000000110011011001101,
    24'b000000110110011011001100,
    24'b000000010110011011000100,
    24'b000000010110010111001111,
    24'b000001000110010111001101,
    24'b000010010110011111001000,
    24'b000010100110011111001001,
    24'b000010100110011011000100,
    24'b000010010110011011000001,
    24'b000010000110010110111110,
    24'b000010010110011011000010,
    24'b000001110110010111000010,
    24'b000001010110001111000101,
    24'b000001100110010111001110,
    24'b000001000110011111001110,
    24'b000000100110100011001101,
    24'b000000010110100011001111,
    24'b000000000110011011010010,
    24'b000000010110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010010,
    24'b000000100110011011010010,
    24'b000000010110011011001111,
    24'b000000010110011011001110,
    24'b000000000110011011010001,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001111,
    24'b000000010110011011001111,
    24'b000000010110011011001111,
    24'b000000010110011111001111,
    24'b000000010110011011010001,
    24'b000000010110011111010000,
    24'b000000100110011011010001,
    24'b000000010110011011010011,
    24'b000000000110011011010010,
    24'b000000000110011111001111,
    24'b000000010110100011001111,
    24'b000000100110011011010100,
    24'b000000010110100011001100,
    24'b000000010110010111001110,
    24'b000000110110011011001111,
    24'b000000110110011111001101,
    24'b000000100110011011010010,
    24'b000000110110100011001110,
    24'b000000110110011111001111,
    24'b000001000110011111001110,
    24'b000000100110010111001101,
    24'b000000100110011111001101,
    24'b000000110110011011010000,
    24'b000000100110100011010000,
    24'b000000010110100011010110,
    24'b000000010110100011001100,
    24'b000000100110011011010001,
    24'b000000110110010111001111,
    24'b000000010110011111001111,
    24'b000000010110011011010010,
    24'b000000000110011011010011,
    24'b000000010110011011010011,
    24'b000000010110011011001111,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011111010100,
    24'b000000000110011011010100,
    24'b000000110110010111010010,
    24'b000000110110010111010000,
    24'b000001000110011011010001,
    24'b000000110110010111010010,
    24'b000000100110011011010100,
    24'b000000010110010111010011,
    24'b000000010110011011001111,
    24'b000000010110011011001101,
    24'b000000000110100011001011,
    24'b000000000110011111001111,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011011010001,
    24'b000000000110011111010010,
    24'b000000010110011111010011,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011011010000,
    24'b000000100110010111010000,
    24'b000000010110011011010010,
    24'b000000010110011111010101,
    24'b000000010110011011010010,
    24'b000000010110011011001111,
    24'b000000010110011111001011,
    24'b000000000110100011001011,
    24'b000000000110011111001111,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000010110100111001111,
    24'b000000100110100111010010,
    24'b000000100110100111010010,
    24'b000000010110011111010011,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000100110100011010100,
    24'b000000000110100111010110,
    24'b000000100110011111010011,
    24'b000000010110011011010000,
    24'b000000010110100011001101,
    24'b000000010110100011001101,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000
};


assign mem_yellow = memory_yellow;

logic [23:0] memory_red [0:4899] = '{
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100011001100,
    24'b000000000110100011001110,
    24'b000000000110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000010110011011010010,
    24'b000000010110011011010000,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011001111,
    24'b000000000110011011001111,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000010110011111010010,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000100110010111001111,
    24'b000000100110010111010000,
    24'b000000100110010111010000,
    24'b000000100110010111010000,
    24'b000000100110010111001111,
    24'b000000010110100011001111,
    24'b000000010110100011001111,
    24'b000000000110011111001100,
    24'b000000010110100011001101,
    24'b000000000110011111001100,
    24'b000000000110011111001100,
    24'b000000000110011111001100,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011001111,
    24'b000000010110100011001111,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110100011010011,
    24'b000000000110100011010011,
    24'b000000010110011111010011,
    24'b000000010110011111010011,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011011010000,
    24'b000000010110011011010010,
    24'b000000000110011111010001,
    24'b000000010110100011010001,
    24'b000000010110100011010000,
    24'b000000010110100011001111,
    24'b000000000110011111001110,
    24'b000000000110011111001101,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000100110100011001110,
    24'b000000010110011011001111,
    24'b000000100110011111010011,
    24'b000000100110011011010100,
    24'b000000100110011011010101,
    24'b000000000110100011010011,
    24'b000000000110100011010010,
    24'b000000000110100011010000,
    24'b000000000110100011010000,
    24'b000000100110100011001111,
    24'b000000100110100011001111,
    24'b000000010110011111010001,
    24'b000000000110011111001101,
    24'b000000000110011111001101,
    24'b000000010110100111010000,
    24'b000000100110100111010011,
    24'b000001010110100111010100,
    24'b000000110110011111010011,
    24'b000000110110011111010100,
    24'b000000010110011111010011,
    24'b000000100110011111010100,
    24'b000000100110011111010100,
    24'b000000100110011111010001,
    24'b000000100110011111010010,
    24'b000000100110011111010010,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001101,
    24'b000000000110011011001011,
    24'b000000000110010111001110,
    24'b000000010110011011010010,
    24'b000000010110010111010100,
    24'b000000000110010011010100,
    24'b000000010110100011001111,
    24'b000000010110011111001110,
    24'b000001000110011111001101,
    24'b000001000110011011001011,
    24'b000001100110010011001010,
    24'b000001100110010011001001,
    24'b000001110110010111001001,
    24'b000001010110010011000101,
    24'b000001100110011011000100,
    24'b000001100110011011000110,
    24'b000001110110011011001001,
    24'b000001010110010111001001,
    24'b000001000110011011001010,
    24'b000001000110011011001101,
    24'b000001000110011011001111,
    24'b000000110110010111010000,
    24'b000000110110010111010001,
    24'b000000100110011111010001,
    24'b000000100110011111010001,
    24'b000001000110011011010001,
    24'b000000100110011111010001,
    24'b000000000110010111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000010110100011010000,
    24'b000000010110011111010000,
    24'b000000000110011111001101,
    24'b000000000110011011001011,
    24'b000000100110010111001111,
    24'b000001110110101011010111,
    24'b000001000110100111010011,
    24'b000001010110010111001101,
    24'b000001100110010111000111,
    24'b000010100110010111000101,
    24'b000011010110001010111111,
    24'b000101000110001110111100,
    24'b000110000110000110111000,
    24'b000101010101110110110010,
    24'b000100110101101010101101,
    24'b000101010101101010101010,
    24'b000101000101100110100111,
    24'b000101000101100110101010,
    24'b000101110101111110110011,
    24'b000100010110010110110111,
    24'b000010010110001110110111,
    24'b000010000110010011000000,
    24'b000010000110010011000011,
    24'b000001010110001111001000,
    24'b000001000110011011001110,
    24'b000001000110011111001011,
    24'b000001000110011111010000,
    24'b000000100110100011010101,
    24'b000000000110011111001110,
    24'b000000100110011111001111,
    24'b000000000110011111010011,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110100111010011,
    24'b000000000110011111001111,
    24'b000000110110010011001011,
    24'b000000000110010111001101,
    24'b000001100110011111010101,
    24'b000000000110010111001010,
    24'b000010110110101111001000,
    24'b000011000110000011000001,
    24'b000100000110100011000010,
    24'b000110010110000110110111,
    24'b000111110101100110011010,
    24'b000101010100001001111010,
    24'b000010000010100101010111,
    24'b000000000001011100111100,
    24'b000000010000110100110000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001000100111000,
    24'b000000010001110001000110,
    24'b000011000011001101100110,
    24'b000101000100111010001011,
    24'b000110110101110110101000,
    24'b000101000110001010110100,
    24'b000011010110010011001010,
    24'b000001010110010111001100,
    24'b000001010110100011001000,
    24'b000010000110100111001111,
    24'b000000110110010111010010,
    24'b000000000110011011010011,
    24'b000000000110011111010001,
    24'b000000000110100011001100,
    24'b000000100110011111001111,
    24'b000000100110011011010001,
    24'b000000010110011011001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011001111,
    24'b000000000110011011010001,
    24'b000000010110011011001111,
    24'b000001010110011011001111,
    24'b000001000110011011010011,
    24'b000001100110011011010010,
    24'b000011010110010011000110,
    24'b001000000101111110110000,
    24'b000111110100110110001110,
    24'b000010010010001001010100,
    24'b000000010000111100110011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001011010000000000000000,
    24'b101010100010101100110101,
    24'b101011110010111100110110,
    24'b101011100011000000110110,
    24'b101011010010111100110101,
    24'b101010010011000100110111,
    24'b101000110011001100111000,
    24'b001011000000000000000001,
    24'b001010010000000000000010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000100001010000110110,
    24'b000100010011100001110100,
    24'b000111100101110010101010,
    24'b000110010110100011001010,
    24'b000010110110010011001000,
    24'b000001010110011111001100,
    24'b000000110110010111001100,
    24'b000001010110011111001100,
    24'b000000010110011011001001,
    24'b000000100110010111001100,
    24'b000000110110010111010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000010110011111001111,
    24'b000001010110011111001111,
    24'b000000000110011111010110,
    24'b000001010110110111011011,
    24'b000010110110000111000011,
    24'b000111000101111010110000,
    24'b000100000011101001111001,
    24'b000000000001001100111011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010001010000001100000011,
    24'b101010000010001100100001,
    24'b110011000010101000101110,
    24'b110100010010100000101010,
    24'b111011010001101100100110,
    24'b111100000001101000100010,
    24'b111011000001110000100010,
    24'b111011100001101100100100,
    24'b111011010001101100100100,
    24'b111011110001101000100011,
    24'b111011100001101100100100,
    24'b111010110001110000100101,
    24'b111010100001111000100000,
    24'b111011100001101100100011,
    24'b110110000010011000101010,
    24'b110010110010101000101111,
    24'b101001100010000100101101,
    24'b001100110000000000000001,
    24'b000000000000000000000000,
    24'b000000000000111100101111,
    24'b000001100010010101011000,
    24'b000100100101001010010011,
    24'b000101000110001010111011,
    24'b000001100110101011001000,
    24'b000000100110011111001010,
    24'b000000010110001011001101,
    24'b000000010110100011010101,
    24'b000001000110101111011000,
    24'b000000100110010011010010,
    24'b000000010110011011010000,
    24'b000000100110011111010001,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010000,
    24'b000000000110011111010000,
    24'b000000010110011011001101,
    24'b000011000110011011001100,
    24'b000011000110011011000111,
    24'b000101110110010110111000,
    24'b000100100011111001111001,
    24'b000000010001001100110010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100011100001111100100010,
    24'b111000110001111100101101,
    24'b111010000001101100100111,
    24'b111011000001101000101000,
    24'b111011010001101100100110,
    24'b111011000001110000100010,
    24'b111011100001101100100011,
    24'b111010110001110000100110,
    24'b111010100001110000100111,
    24'b111010100001110000100110,
    24'b111010100001110100100100,
    24'b111011000001101100100100,
    24'b111011100001101100100100,
    24'b111011010001101100100101,
    24'b111100000001100100100111,
    24'b111011010001101000100110,
    24'b111011000001110000100011,
    24'b111011010001101000100100,
    24'b111011010001101000100110,
    24'b111010010001111000101001,
    24'b110100110010011000110001,
    24'b100011000010001000100111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000010010010010101010101,
    24'b000101010101011010100000,
    24'b000011010110100011000001,
    24'b000001100110110111010011,
    24'b000001000110010011010001,
    24'b000010000110001011001011,
    24'b000001110110010111001000,
    24'b000000110110011011001110,
    24'b000000110110010111010000,
    24'b000000010110011011010000,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000010110100011010001,
    24'b000000010110100011010001,
    24'b000001000110011011001101,
    24'b000101000110001111000101,
    24'b000101110100111010010100,
    24'b000000000001010000110100,
    24'b000000000000000000000000,
    24'b001010110000000000000010,
    24'b101001010010010100101101,
    24'b111001000001111000100110,
    24'b111011110001101000100011,
    24'b111011000001110000100101,
    24'b111011000001110100100001,
    24'b111011000001110000100100,
    24'b111010110001110000100101,
    24'b111011110001101000100100,
    24'b111011110001101100100011,
    24'b111010110001110100100011,
    24'b111100000001101000100011,
    24'b111011100001101100100011,
    24'b111011000001101100100011,
    24'b111011010001101100100011,
    24'b111011100001101100100011,
    24'b111011010001110000100011,
    24'b111011100001110000100001,
    24'b111011100001101100100100,
    24'b111010100001110000100111,
    24'b111011100001101100100010,
    24'b111011010001110100100001,
    24'b111011100001110000100011,
    24'b111011010001110100100101,
    24'b111011000001111100100101,
    24'b111000000010000000100111,
    24'b100000100001010100011010,
    24'b000000000000000000000000,
    24'b000000100000110000101001,
    24'b000010110011010001100111,
    24'b000110010110000110110011,
    24'b000011010110010111001011,
    24'b000001010110010011010000,
    24'b000000100110100011010010,
    24'b000000110110011011001110,
    24'b000000110110011011001110,
    24'b000000010110011011010000,
    24'b000000100110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011010000,
    24'b000000000110011011010011,
    24'b000000100110011011010100,
    24'b000000010110011011001110,
    24'b000000000110100011010101,
    24'b000000100110100011010110,
    24'b000010000110010111010000,
    24'b000001110110100011001111,
    24'b000101100110001110110011,
    24'b000100000011001101101101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101111010010101000110101,
    24'b111000110001111100100111,
    24'b111010110001110000100101,
    24'b111011000001101100100101,
    24'b111011000001101100100100,
    24'b111011010001101100100100,
    24'b111011010001110000100011,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011000001110000100011,
    24'b111011100001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011100001101100100100,
    24'b111011010001101100100101,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b110111100010000100101011,
    24'b011101000001101000011111,
    24'b000000000000000000000000,
    24'b000000100001011100111100,
    24'b000110100101100010100100,
    24'b000010000110010111000110,
    24'b000001100110100011001110,
    24'b000001000110101011010101,
    24'b000000000110011011010100,
    24'b000000010110011111010001,
    24'b000000100110100111001111,
    24'b000000000110010111001110,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011010000,
    24'b000000000110011011010011,
    24'b000000000110011011001111,
    24'b000000100110011011001110,
    24'b000000110110011011001100,
    24'b000000000110100011001111,
    24'b000001110110010111000010,
    24'b000101110101111010100110,
    24'b000000100010001101010010,
    24'b000000000000000000000000,
    24'b010100010000110000010010,
    24'b110110010010000000101100,
    24'b111100000001101100100010,
    24'b111010110001110000100011,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010110001111100100110,
    24'b110011110010011100110101,
    24'b001010000000011000010001,
    24'b000000000000111000101001,
    24'b000110000100010101111101,
    24'b000101110110011010111100,
    24'b000001000110100011001110,
    24'b000001000110011011001101,
    24'b000001100110010111001101,
    24'b000001000110100111001110,
    24'b000000000110011011001111,
    24'b000000100110010111010001,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000100110011111010001,
    24'b000000110110011011001110,
    24'b000000010110011011010000,
    24'b000000010110011111001100,
    24'b000001100110000010111101,
    24'b000101000101011110011100,
    24'b000000100001011100111110,
    24'b000000000000000000000000,
    24'b011110000001010100011000,
    24'b111010100001111000101001,
    24'b111011110001110000100101,
    24'b111101000001111000101000,
    24'b111011010001110000100001,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101000100001,
    24'b111001100001111100100101,
    24'b111000110010000100101001,
    24'b010011010000001100000100,
    24'b000000000000000000000000,
    24'b000010000011100101110001,
    24'b000011010110010110111010,
    24'b000010110110001111001010,
    24'b000000110110001111010000,
    24'b000000000110101111010010,
    24'b000000000110011111001110,
    24'b000000010110011011010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010011,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110010111001111,
    24'b000000010110010111010000,
    24'b000000100110011111010001,
    24'b000000000110011111010010,
    24'b000000010110100011010001,
    24'b000010100110010111001100,
    24'b001001000101011010100100,
    24'b000000000000101100101101,
    24'b000000000000000000000000,
    24'b101111100010110000110011,
    24'b111010100001111000101001,
    24'b111001110001101100100011,
    24'b111010110001101100101000,
    24'b111010110001110000100100,
    24'b111011010001101100100110,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100101,
    24'b111011010001101100101000,
    24'b111010110001110000100011,
    24'b111001000001111100011111,
    24'b100100110010001100101100,
    24'b000000000000000000000000,
    24'b000110000011101101110101,
    24'b000101000110001010111100,
    24'b000001000110011111011000,
    24'b000001000110100111010101,
    24'b000000110110011011001100,
    24'b000000110110011011010000,
    24'b000000000110011111001110,
    24'b000000010110100011001111,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110010111010001,
    24'b000000110110100011010010,
    24'b000001000110011111001110,
    24'b000001000110011011001101,
    24'b000010100110010111000011,
    24'b000111100101110110101010,
    24'b000000010001010100111010,
    24'b000000000000000000000000,
    24'b101111100010011100110111,
    24'b111011110001100100100000,
    24'b111011000001100100100101,
    24'b111011100001101100100100,
    24'b111010010001110100100010,
    24'b111011110001101000100011,
    24'b111010110001110000100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010110001110000100011,
    24'b111101000001011100100110,
    24'b111011010001101100100010,
    24'b111011110001101100100100,
    24'b111010110001110000100111,
    24'b100111010010010000100110,
    24'b000000000000000000000000,
    24'b000011000011110101101111,
    24'b000100010110010010111101,
    24'b000001110110010111001110,
    24'b000001010110010111010000,
    24'b000000000110100011010001,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010011,
    24'b000000100110011011001111,
    24'b000001010110011111001111,
    24'b000001100110011011000110,
    24'b000101100110001110101111,
    24'b000000100001001001000000,
    24'b000000000000000000000000,
    24'b101111010010011000110000,
    24'b111011000001110000100010,
    24'b111010100001110000100110,
    24'b111011010001101000100001,
    24'b111011010001101000100100,
    24'b111011100001101000100110,
    24'b111011000001110000100011,
    24'b111011010001101100100011,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010100001110000100111,
    24'b111011100001101100100100,
    24'b111011000001110000100101,
    24'b111010110001110000100010,
    24'b111010100001110000101001,
    24'b111001100001110000100110,
    24'b100110000001110100101010,
    24'b000000000000000000000000,
    24'b000110110100110010001001,
    24'b000100000110000011000100,
    24'b000000010110011011010001,
    24'b000000100110010111010000,
    24'b000000010110011111010101,
    24'b000000000110011011010010,
    24'b000000000110011111010001,
    24'b000000000110011111001110,
    24'b000000000110011111001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010010,
    24'b000000010110011011001111,
    24'b000000110110011011001101,
    24'b000000000110100011010100,
    24'b000001110110100111010000,
    24'b000001100110010011001000,
    24'b000101000110010010111110,
    24'b000001110010101001011100,
    24'b000000000000000000000000,
    24'b101100000011000000110111,
    24'b111011010001101100011111,
    24'b111011010001101000100111,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111001110010000000100110,
    24'b010011100000101000001011,
    24'b000000110000110100101111,
    24'b000110110101101110100001,
    24'b000010010110101011001001,
    24'b000001100110100011001110,
    24'b000001100110011111010101,
    24'b000000010110010111010101,
    24'b000000010110011011010011,
    24'b000000010110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001100,
    24'b000000000110100011001011,
    24'b000000010110011111010000,
    24'b000000000110001111001011,
    24'b000011000110001010111000,
    24'b000011010100010001111001,
    24'b000000000000000000000000,
    24'b011100010001000100010110,
    24'b111001000001111000100010,
    24'b111011000001101100100100,
    24'b111010010001111000100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011110001100100011111,
    24'b110111010010001000101111,
    24'b001100100000011100001010,
    24'b000000000001110000111110,
    24'b000110100110000110110011,
    24'b000011100110010111001011,
    24'b000000100110001111010001,
    24'b000001000110011011010001,
    24'b000000110110010111010000,
    24'b000000100110010111010010,
    24'b000000010110011111010101,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010000,
    24'b000000010110011111010011,
    24'b000000010110011111010000,
    24'b000000110110011111010011,
    24'b000010010110010011001100,
    24'b000110010101101010100011,
    24'b000000010000111100101011,
    24'b000000000000000000000000,
    24'b111000100010001000100110,
    24'b111010110001110100100101,
    24'b111011010001101000100101,
    24'b111011110001110000100011,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010100001110000100001,
    24'b111011000001100100100011,
    24'b110010010010110000101110,
    24'b000000000000000000000000,
    24'b000010110011001101101000,
    24'b000011010101111011000001,
    24'b000001100110100111010110,
    24'b000000000110011111010000,
    24'b000000110110011011001110,
    24'b000001000110010111001111,
    24'b000000010110011111010011,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110010111010100,
    24'b000000010110010111010101,
    24'b000001000110001111010001,
    24'b000101100110000110111100,
    24'b000001110010100101011111,
    24'b000000000000000000000000,
    24'b110000110010110000110011,
    24'b111010100001100000100001,
    24'b111011010001101100100110,
    24'b111010010001110100100101,
    24'b111011010001101100100010,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011100001101000101000,
    24'b111100000001101000100101,
    24'b111010110001110100100011,
    24'b100000100001101000011111,
    24'b000000000000000000000000,
    24'b000110000101101010100011,
    24'b000010010110011111001001,
    24'b000000000110011111010100,
    24'b000000010110011111010000,
    24'b000001000110011011001011,
    24'b000000010110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000110110011011001100,
    24'b000001010110001111010100,
    24'b000001100110001111001010,
    24'b000111000101011010010111,
    24'b000000010000111000101001,
    24'b010110000001010000010110,
    24'b111011100001011100100101,
    24'b111100000001101000100100,
    24'b111011100001101000100110,
    24'b111010110001110000100010,
    24'b111010110001110000100101,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010110001110000100110,
    24'b111010110001110000100101,
    24'b111011000001101100100101,
    24'b110111000001111100101000,
    24'b000000000000000000000000,
    24'b000001000010010001001000,
    24'b000110010110011110111000,
    24'b000001010110010111010100,
    24'b000000010110100011010010,
    24'b000000110110011111001001,
    24'b000000000110011111010010,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000010110011111001111,
    24'b000000100110011111010011,
    24'b000000000110011111010010,
    24'b000000110110100011001100,
    24'b000000100110000111001101,
    24'b000100100110010010111110,
    24'b000001100010010001001101,
    24'b000000000000000000000000,
    24'b110100010010011100101110,
    24'b111011000001101000100110,
    24'b111010100001110000100100,
    24'b111011000001101100100100,
    24'b111011010001110000100010,
    24'b111011010001101100100110,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011110001101000100010,
    24'b111010100001110100100100,
    24'b111100000001100100100111,
    24'b111011010001101100100011,
    24'b100101110001110000100110,
    24'b000000000000000000000000,
    24'b001001000101111110011111,
    24'b000001110110011011001011,
    24'b000001010110011111010010,
    24'b000000100110100111010011,
    24'b000000010110100011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000010110011111001101,
    24'b000000100110011011010011,
    24'b000000100110010111010010,
    24'b000000100110011111001000,
    24'b000100000110110111010001,
    24'b001000010101101010100011,
    24'b000000000000000000000000,
    24'b010101100001001000010101,
    24'b111001010001111000100111,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100110,
    24'b111010100001110100100010,
    24'b111011110001100100101000,
    24'b111011010001110000100001,
    24'b110110100010010000101110,
    24'b000000000000000000000000,
    24'b000000010010011001010101,
    24'b000110100110110111000100,
    24'b000010110110001011001111,
    24'b000000000110011111010011,
    24'b000000010110011111001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111001111,
    24'b000000010110011011010010,
    24'b000001000110010011010000,
    24'b000000100110100111000101,
    24'b000011000110000110111011,
    24'b000011000010100101011011,
    24'b000000000000000000000000,
    24'b110011000010100100110000,
    24'b111011100001101100100011,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010110001101100101001,
    24'b111011100001101100100001,
    24'b111011100001101100100100,
    24'b111011000001110000100000,
    24'b111011100001101100100001,
    24'b100111000010011000101100,
    24'b000000000000000000000000,
    24'b001000110110000010101100,
    24'b000010110110010111001111,
    24'b000001010110010011001111,
    24'b000000000110011111001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000110110010111001110,
    24'b000000000110101111001000,
    24'b000110110110011010110111,
    24'b000000000000100000101001,
    24'b000000000000000000000000,
    24'b111010100001110100100101,
    24'b111011010001101100100011,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010110001101100100111,
    24'b111011010001101100100001,
    24'b111011000001101100100101,
    24'b111011010001101100100110,
    24'b111011100001101100100011,
    24'b110101100010010100101111,
    24'b000000000000000000000000,
    24'b000111100100100110000110,
    24'b000010000110010111000111,
    24'b000001100110010011010001,
    24'b000000000110011111010010,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110010111010100,
    24'b000000010110011011010001,
    24'b000000110110011011001110,
    24'b000001000110100011001100,
    24'b000110100101011110010111,
    24'b000000000000000000000000,
    24'b100100100010000100100100,
    24'b111011000001111100100110,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010110001110000100010,
    24'b111011010001101100100100,
    24'b111010110001110000100110,
    24'b111011010001101100100101,
    24'b111010100001110000100110,
    24'b111010100001110000101000,
    24'b001011110000000000000001,
    24'b000000000001011101000101,
    24'b000101000110010110111011,
    24'b000001000110011011010001,
    24'b000000010110011111010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011011010001,
    24'b000000000110010111010101,
    24'b000000010110011011010000,
    24'b000000100110011011001010,
    24'b000100000110010011001000,
    24'b000000110010110001011100,
    24'b000000000000000000000000,
    24'b110110010010001100101010,
    24'b111011100001100100100011,
    24'b111011010001101100100101,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010110001110100100001,
    24'b111011100001101000100111,
    24'b111010100001110000100101,
    24'b111011010001110000100001,
    24'b111011010001101100100010,
    24'b111011110001101000100011,
    24'b101010010011001100111110,
    24'b000000010001000000110100,
    24'b000110010110000010101000,
    24'b000010000110010011001100,
    24'b000000000110011111001101,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110011011010001,
    24'b000000010110011011010000,
    24'b000000010110011011001101,
    24'b000011110110000110111100,
    24'b000000010001001100110010,
    24'b000000000000000000000000,
    24'b111000010010001000101000,
    24'b111011110001100100100110,
    24'b111011010001101100100101,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010110001110000100100,
    24'b110101110010001100101001,
    24'b000000000000000000000000,
    24'b000111100101010110010011,
    24'b000010100110010111000111,
    24'b000000000110011011010100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000110110011011001011,
    24'b000101000101110010101110,
    24'b000000000000000000000000,
    24'b010000010000000000000001,
    24'b111010110001111100101000,
    24'b111011100001101100100010,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101000100100,
    24'b111010010001110100101010,
    24'b000000000000000000000000,
    24'b000100000011101101110011,
    24'b000010010110100011000011,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000001000110010111001011,
    24'b001000110101111110100101,
    24'b000000000000000000000000,
    24'b101001010010000100101001,
    24'b111011000001101000100110,
    24'b111010110001110000100001,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011000001110000100101,
    24'b001111010000010000000100,
    24'b000000000001111101001110,
    24'b000010000110011110111100,
    24'b000000110110011011001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110010111001111,
    24'b000000010110011011010000,
    24'b000001010110010111001010,
    24'b001001110101000010010000,
    24'b000000000000000000000000,
    24'b101001110010001000100110,
    24'b111011010001101000101000,
    24'b111010110001110000100100,
    24'b111011000001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100011,
    24'b111011100001101100100100,
    24'b010100100000001100000011,
    24'b000000000001001000111000,
    24'b000100110110000010110111,
    24'b000000110110011011001110,
    24'b000000000110011111010001,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011011001111,
    24'b000000000110010111010000,
    24'b000001110110011011001010,
    24'b000110010011110101110100,
    24'b000000000000000000000000,
    24'b110011000010100000110010,
    24'b111011100001101000100110,
    24'b111011010001101100100011,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011000001101100100100,
    24'b111010000001111000100111,
    24'b110010000010101000110110,
    24'b000000000000111000101100,
    24'b000101000110000110111000,
    24'b000001000110011011001110,
    24'b000000000110011011010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000010110011111001111,
    24'b000000010110011011001111,
    24'b000010010110011011001000,
    24'b000011110011001001100101,
    24'b000000000000000000000000,
    24'b110100010010011000101111,
    24'b111010110001110000100101,
    24'b111011100001101100100011,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111100000001110000100111,
    24'b110011100010010100110001,
    24'b000000000000101100101000,
    24'b000101110110000110110100,
    24'b000000110110010111001110,
    24'b000000010110011011010001,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000010110011111001111,
    24'b000001010110100011010000,
    24'b000011000110011011001010,
    24'b000010000010110001011110,
    24'b000000000000000000000000,
    24'b110100010010011100101101,
    24'b111011010001101100100110,
    24'b111011010001101000100101,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100011,
    24'b110010000010101100110011,
    24'b000000000000000000000000,
    24'b000101110110000110101101,
    24'b000001000110010011001111,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010000,
    24'b000001010110011111010010,
    24'b000011010110011011001011,
    24'b000001110010100101011010,
    24'b000000000000000000000000,
    24'b110100000010100000101100,
    24'b111011100001101100100100,
    24'b111011010001101100100011,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010110001110000100010,
    24'b110001100010110000110011,
    24'b000000000000000000000000,
    24'b000110010101111110101101,
    24'b000000100110011011001101,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000010110011111010010,
    24'b000001010110011111010011,
    24'b000011000110011011001011,
    24'b000001010010111001011110,
    24'b000000000000000000000000,
    24'b110101010010011000101100,
    24'b111011010001110000100010,
    24'b111011010001101100100011,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011100001110100100010,
    24'b110011110010011000110110,
    24'b000000000000011000101010,
    24'b000101100101111110101111,
    24'b000000010110011111001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010001,
    24'b000001000110011011010010,
    24'b000010100110011011001010,
    24'b000010110011110001101100,
    24'b000000000000000000000000,
    24'b110011100010100100110000,
    24'b111011010001110000100010,
    24'b111011010001101100100100,
    24'b111011100001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011100001101100100100,
    24'b111011010001111000100100,
    24'b110001000010101000111010,
    24'b000000000000101100110010,
    24'b000100110110001010110011,
    24'b000000010110100011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010011,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000010110011111001111,
    24'b000001010110100011010000,
    24'b000010000110011011001000,
    24'b001000010100111110000110,
    24'b000000000000000000000000,
    24'b101010010010001000100101,
    24'b111100000001101000100100,
    24'b111011000001110000100110,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011100001101000100100,
    24'b111001110001110100100101,
    24'b010100000000001100000011,
    24'b000000000000110100111001,
    24'b000100100110001110111000,
    24'b000000010110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111001111,
    24'b000000010110011111001100,
    24'b000000010110010111000111,
    24'b000111110101100010011011,
    24'b000000000000000000000000,
    24'b101000110010010100101011,
    24'b111100110001100100100101,
    24'b111011000001110100100010,
    24'b111011010001101100100011,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011000001101100100100,
    24'b111010010001110000100110,
    24'b010001110000001100000100,
    24'b000000000001010101000011,
    24'b000011010110001010111011,
    24'b000000010110011011001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011111001111,
    24'b000000100110011111001101,
    24'b000000100110010111001011,
    24'b000111110101110110101011,
    24'b000000000000000000000000,
    24'b010001010000000000000000,
    24'b111010000001111000100110,
    24'b111011000001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010110001110000100100,
    24'b111010000001111000100111,
    24'b000000000000000000000000,
    24'b000010110011001001100011,
    24'b000010110110001011000100,
    24'b000000100110011011001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000100110011111001111,
    24'b000000110110010111001111,
    24'b000110000101111110110011,
    24'b000000000000111100110001,
    24'b000000000000000000000000,
    24'b111001010001111100100101,
    24'b111010110001100100100110,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010010001100100101011,
    24'b000000000000000000000000,
    24'b000111010100111110001011,
    24'b000010100110001011001001,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011001111,
    24'b000000000110011111001110,
    24'b000000100110011111001111,
    24'b000000000110010111001101,
    24'b000100000110001010110111,
    24'b000000100001111001001011,
    24'b000000000000000000000000,
    24'b110111010001111100101010,
    24'b111011100001110100100011,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101000100100,
    24'b101010100011000000110110,
    24'b000000000000000000000000,
    24'b001000100101011110100110,
    24'b000010000110011111001010,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111001110,
    24'b000000010110100011001101,
    24'b000000000110011011001101,
    24'b000000010110010111001111,
    24'b000000110110100111010010,
    24'b000010100110100011000011,
    24'b000101110100101110000111,
    24'b000000000000000000000000,
    24'b100011100001111000100101,
    24'b111011010001111000100010,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101000100110,
    24'b001101000000000000000001,
    24'b000000000000110100110100,
    24'b000110010110001110111111,
    24'b000001010110011111001100,
    24'b000000010110010011001110,
    24'b000000010110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111001110,
    24'b000000000110011111001100,
    24'b000000000110011011001101,
    24'b000000000110010011001110,
    24'b000001110110100111010100,
    24'b000001010110010111001011,
    24'b000111100110001110110000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111010010001110100100110,
    24'b111011000001110000100011,
    24'b111011100001101100100011,
    24'b111011010001101100100101,
    24'b111011100001101100100011,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011000001110000100100,
    24'b111011000001101100100011,
    24'b111011100001101000100101,
    24'b110100110010011100101011,
    24'b000000000000000000000000,
    24'b000011110010100101100101,
    24'b000011110110001111000101,
    24'b000000110110100111010110,
    24'b000000000110100011001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000001100110100111010010,
    24'b000000110110011111010101,
    24'b000101010110100011000001,
    24'b000000110001110101001011,
    24'b000000000000000000000000,
    24'b110010010010110000110001,
    24'b111011000001110100100010,
    24'b111011110001101000100101,
    24'b111011000001101100100111,
    24'b111011110001101100100011,
    24'b111010110001110000100101,
    24'b111011110001101000100110,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011100001101100100101,
    24'b111011100001101100100100,
    24'b111010100001110100100101,
    24'b111010100001101100100000,
    24'b111011010001100100100111,
    24'b100111110010011000101000,
    24'b000000000000000000000000,
    24'b000111000100111110011100,
    24'b000010010110001111001010,
    24'b000000110110011111010011,
    24'b000000100110011111010001,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000100110011111010001,
    24'b000000010110100011010101,
    24'b000001010110010011010010,
    24'b000011100110001111000111,
    24'b000110010100100110001001,
    24'b000000000000000000000000,
    24'b010110010001001000010100,
    24'b111010100001110100100101,
    24'b111010110001101100101000,
    24'b111010110001110000100011,
    24'b111011010001101000101001,
    24'b111010000001111000100010,
    24'b111011110001101000100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010100001110000100010,
    24'b111100010001100100100101,
    24'b111100000001100100100100,
    24'b111011000001101100100110,
    24'b111000000001111100100111,
    24'b000000000000000000000000,
    24'b000000010001100100111111,
    24'b000111000110110111000010,
    24'b000000110110001111001001,
    24'b000000100110011011010001,
    24'b000000100110011011010010,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000100110011111010001,
    24'b000000100110100011010010,
    24'b000000000110011011010010,
    24'b000001110110001111010000,
    24'b000001000110011011000111,
    24'b000111000110010010110011,
    24'b000000110001010100111101,
    24'b000000000000000000000000,
    24'b110100010010011100110000,
    24'b111010110001110000100001,
    24'b111011100001101000100001,
    24'b111011100001101000100111,
    24'b111011010001110000100010,
    24'b111010110001110000100110,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010110001110000100010,
    24'b111010100001110100100011,
    24'b111100000001101000100111,
    24'b111010110001111100100100,
    24'b100101000001111100100010,
    24'b000000000000000000000000,
    24'b000100010100101110000111,
    24'b000001010110100111001000,
    24'b000000100110010111001000,
    24'b000000110110011111001110,
    24'b000000010110010111010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000100110011011010000,
    24'b000000110110100011010100,
    24'b000001010110011011001000,
    24'b000011110110010010111111,
    24'b000011100011110001111011,
    24'b000000000000000000000000,
    24'b010101010001010000010100,
    24'b111100000001101000100001,
    24'b111011010001101100100010,
    24'b111011010001110000100010,
    24'b111011010001101100100100,
    24'b111011100001101000100110,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011100001101100100100,
    24'b111011000001110000100001,
    24'b111100010001011100101010,
    24'b110111100010001000101000,
    24'b000000000000000000000000,
    24'b000000010000111000110110,
    24'b000111100110010110110100,
    24'b000001000110101111010010,
    24'b000000110110011011001011,
    24'b000000100110100011001011,
    24'b000000000110100011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010001,
    24'b000000100110100011010111,
    24'b000000110110010111010010,
    24'b000010000110011011001001,
    24'b000110100110010110111000,
    24'b000000000001011001000010,
    24'b000000000000000000000000,
    24'b110000100010101000110011,
    24'b111001110001101100100100,
    24'b111011010001101100101000,
    24'b111011110001101100100001,
    24'b111010110001110000100110,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010110001110000100100,
    24'b111011000001101100101000,
    24'b100001000001101000011111,
    24'b000000000000000000000000,
    24'b000101010100100010001100,
    24'b000011100110001111000000,
    24'b000000000110010011010011,
    24'b000000010110011011001111,
    24'b000000110110011011001011,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110010011011000,
    24'b000000100110011011011010,
    24'b000001000110101111010010,
    24'b000100010110101011000100,
    24'b000101110100101010010000,
    24'b000000000000000000000000,
    24'b001010100000001000001010,
    24'b111000010010000100101100,
    24'b111010100001110000100101,
    24'b111011000001110000100101,
    24'b111010100001110100100010,
    24'b111011000001110000100010,
    24'b111011110001101000100010,
    24'b111011000001110000100010,
    24'b111100000001101000100010,
    24'b111010110001110000100100,
    24'b111011100001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010100001110000100101,
    24'b111011010001101000100101,
    24'b111011010001101100100011,
    24'b111010110001110000100010,
    24'b111010100001110100100011,
    24'b111011100001101000100101,
    24'b111010000001110100100100,
    24'b111100010001101000100010,
    24'b110001110010101100110000,
    24'b000000000000000000000000,
    24'b000000110001100001001010,
    24'b000101010110001010111100,
    24'b000001100110011011001100,
    24'b000000100110011011010011,
    24'b000000010110011011010010,
    24'b000000010110011011001111,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010001,
    24'b000000100110010111010100,
    24'b000000000110011111010001,
    24'b000001100110010011000100,
    24'b000110110110001010111101,
    24'b000010010010100101011001,
    24'b000000000000000000000000,
    24'b011111010001001000011000,
    24'b111000000010000100100011,
    24'b111100100001100100100101,
    24'b111100100001100100100111,
    24'b111011010001101100100101,
    24'b111011010001101100100110,
    24'b111010010001110100100101,
    24'b111011010001101100100011,
    24'b111011100001101100100100,
    24'b111011000001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011100001101000100101,
    24'b111011000001110000100100,
    24'b111011110001101000100100,
    24'b111011110001101000100110,
    24'b111101000001101000101000,
    24'b111010010001111100101001,
    24'b001101010000100000001010,
    24'b000000000000110100101010,
    24'b000110000101011110011111,
    24'b000010000110100011001001,
    24'b000001100110101111010101,
    24'b000000000110010111001111,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001101,
    24'b000000110110011011001100,
    24'b000001000110010011010010,
    24'b000000000110001011010001,
    24'b000001000110011111010001,
    24'b000011110110010011001101,
    24'b000111000101100110101110,
    24'b000000000001010000111000,
    24'b000000000000000000000000,
    24'b101011110010111100111000,
    24'b111011100001110000100000,
    24'b111010110001110100100101,
    24'b111011100001101100100101,
    24'b111011010001101100100110,
    24'b111011000001101100100111,
    24'b111011100001101000100110,
    24'b111011010001110000100010,
    24'b111011100001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001110000100001,
    24'b111011100001101100100011,
    24'b111011010001101100101000,
    24'b111011100001101000100101,
    24'b111011000001110000100010,
    24'b111011000001110000100011,
    24'b111010000010000100101001,
    24'b100000000001111100100100,
    24'b000000000000000000000000,
    24'b000101110100000001111111,
    24'b000011010110011011000101,
    24'b000000010110011111001101,
    24'b000000100110011111010001,
    24'b000000100110011111010001,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000010110011011010011,
    24'b000001000110010011010101,
    24'b000000010110011011010100,
    24'b000000000110011011001111,
    24'b000010000110100111001110,
    24'b000001110110100011000110,
    24'b000101110101001110010010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110000010010100000101101,
    24'b111010100001111000100110,
    24'b111010000001111000100001,
    24'b111100100001101100100001,
    24'b111010010001111100100101,
    24'b111011100001101000101000,
    24'b111010010001110100100100,
    24'b111011000001101100100011,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010110001110000100010,
    24'b111011000001110000100101,
    24'b111011100001101000100111,
    24'b111010100001110000100001,
    24'b111011010001110000100010,
    24'b111010000001110100101000,
    24'b100101010010000100100011,
    24'b000000000000000000000000,
    24'b000010010010011001011011,
    24'b000110000110000010110101,
    24'b000000100110010111001100,
    24'b000000110110011111010100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110010111010101,
    24'b000000010110010111010100,
    24'b000000010110011111010001,
    24'b000000000110011011001100,
    24'b000001000110011011001011,
    24'b000010000110011111000101,
    24'b000100100110001111000110,
    24'b000110010011111110000101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110000010010011000110001,
    24'b111010110001100000100101,
    24'b111011100001110000100000,
    24'b111011100001101000100000,
    24'b111011100001101000100110,
    24'b111011010001101100100100,
    24'b111011100001101100100011,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010100001110100100010,
    24'b111011110001101000100110,
    24'b111011000001101100100101,
    24'b111011010001110000100001,
    24'b111001110001101100101011,
    24'b100101010010010000101101,
    24'b000000000000000000000000,
    24'b000000100001101001000101,
    24'b000100110110010010101111,
    24'b000001110110011011001001,
    24'b000000010110100011000111,
    24'b000000010110010111010011,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100011001110,
    24'b000000000110100111001101,
    24'b000000010110011011001110,
    24'b000000110110011011010001,
    24'b000001100110001111010010,
    24'b000001010110001011001111,
    24'b000000100110100111010000,
    24'b000011000110001111000001,
    24'b000110000100000101111110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101111110010101100110001,
    24'b111011000001101100100111,
    24'b111011010010000000100100,
    24'b111010110001110000100110,
    24'b111011100001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011100001101100100010,
    24'b111011110001101000100100,
    24'b111011000001110000100011,
    24'b111001110001110100100100,
    24'b100101000010001100101000,
    24'b000000000000000000000000,
    24'b000000010001011101000000,
    24'b000110110101101110101010,
    24'b000001100110010111000011,
    24'b000001100110101011010010,
    24'b000000010110011111010111,
    24'b000000010110100011001000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011111010101,
    24'b000000010110011111010101,
    24'b000001000110011111001011,
    24'b000000110110010011001100,
    24'b000001100110010111001111,
    24'b000100110110001010111111,
    24'b000100100011111101111010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b011111100001010000010110,
    24'b111001110010000000101010,
    24'b111010110001100000011111,
    24'b111011010001111000100110,
    24'b111011100001101100100100,
    24'b111011010001101000100111,
    24'b111011100001101000101000,
    24'b111011010001101100100101,
    24'b111011010001110000100010,
    24'b111100000001101000100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011000001101100100100,
    24'b111011010001101100100100,
    24'b111010100001110000100110,
    24'b111011000001101100100110,
    24'b111011010001101100100110,
    24'b111010010001110100100110,
    24'b111011000001101100100100,
    24'b111011100001101000100110,
    24'b111100000001101000100110,
    24'b111011100001101100100100,
    24'b111011100001101100100010,
    24'b111011100001101100101000,
    24'b111011100001101100100010,
    24'b111000000001111100101011,
    24'b010011000000010000000100,
    24'b000000000000000000000000,
    24'b000000010001101001000000,
    24'b000011100110000110110000,
    24'b000010010110001110111111,
    24'b000000110110010111001010,
    24'b000000000110011011001110,
    24'b000000010110100011001110,
    24'b000000000110011111001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000110110100011010100,
    24'b000000010110010111010001,
    24'b000000000110011011010011,
    24'b000010100110101011010001,
    24'b000101100110000010110110,
    24'b000101010100011110001001,
    24'b000000000000110100110000,
    24'b000000000000000000000000,
    24'b010100010000110000001100,
    24'b110111100010001000101110,
    24'b111010100001101000100101,
    24'b111011100001101100100011,
    24'b111010110001110100100001,
    24'b111011010001110000011111,
    24'b111011100001101100100010,
    24'b111010010001110100100100,
    24'b111011000001110000100011,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011000001101100100100,
    24'b111011110001101000100100,
    24'b111011000001101100100100,
    24'b111100000001101000100100,
    24'b111011010001101100100100,
    24'b111100010001100100100100,
    24'b111100010001101000100011,
    24'b111011000001110100100000,
    24'b111010010001110100100101,
    24'b111011000001101100100111,
    24'b111010110001110000100011,
    24'b111010110001101000011110,
    24'b110010010010110000110100,
    24'b001010110000011000001010,
    24'b000000000000000000000000,
    24'b000000100010001001000111,
    24'b000100110101110110101011,
    24'b000010110110010011000100,
    24'b000010010110100011001110,
    24'b000000010110010111010011,
    24'b000000000110011111010111,
    24'b000000000110011011010100,
    24'b000000010110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000010110100011001111,
    24'b000000000110011111001110,
    24'b000000010110011111010101,
    24'b000000110110100011010100,
    24'b000000000110011011001110,
    24'b000000010110100011010010,
    24'b000001010110010111001101,
    24'b000011110110010011000111,
    24'b000101110101001010010011,
    24'b000000110001001100111010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101111100010110000110100,
    24'b111000110001111100100110,
    24'b111010110001101100100111,
    24'b111011010001101100101000,
    24'b111010110001110000100100,
    24'b111011110001101000100011,
    24'b111011100001101000100110,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010010001110000100110,
    24'b111011110001101000100100,
    24'b111001010001111100100010,
    24'b111011100001101100100010,
    24'b111011000001110000100010,
    24'b111011000001110000100100,
    24'b111010010001110100100101,
    24'b111011100001101100100101,
    24'b111011110001101100011110,
    24'b111011100001101100100010,
    24'b110111100010000100101100,
    24'b011110000001100000011010,
    24'b000000000000000000000000,
    24'b000000100000100000101010,
    24'b000011000011010001101001,
    24'b000111000110011110110000,
    24'b000001110110101111001111,
    24'b000000110110011011001110,
    24'b000000010110010111010001,
    24'b000000000110011111010101,
    24'b000000010110101011011001,
    24'b000000000110010111010011,
    24'b000000000110010111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000010110100011010010,
    24'b000000010110011111001110,
    24'b000000010110100011001011,
    24'b000000010110100011001011,
    24'b000000110110011011001101,
    24'b000001000110010111001111,
    24'b000001100110011011000101,
    24'b000111100110001010101101,
    24'b000010010010100101010110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001101100000000000000001,
    24'b101011110010011000101110,
    24'b111001000010000100100110,
    24'b111011000001110000100011,
    24'b111011110001100100100101,
    24'b111010010001110100100000,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011000001101100100110,
    24'b111100000001101000100100,
    24'b111011110001101100100010,
    24'b111011100001111000100100,
    24'b111011000001111100100110,
    24'b111100000001100100100101,
    24'b111011010001101100100011,
    24'b111010110001110000100100,
    24'b111000100001111100101100,
    24'b100001010001010100010110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001011000111011,
    24'b000101000100110010010011,
    24'b000001100110100010111100,
    24'b000000010110011011001000,
    24'b000000100110011011010011,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000010110011011001111,
    24'b000000110110011011001101,
    24'b000000010110011011001101,
    24'b000000010110011111001100,
    24'b000000100110001111001110,
    24'b000010010110011011001010,
    24'b000100100110010110111010,
    24'b000110100100110110010100,
    24'b000000010001010001000101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001011110000000000000001,
    24'b101011100010000100100110,
    24'b111000110001111100101000,
    24'b111011100001101100100111,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111011000001101100100110,
    24'b111010110001110000100100,
    24'b111011010001110000100010,
    24'b111010000001110000100011,
    24'b111100000001011100100110,
    24'b111001010010000000101000,
    24'b111000110001111100101001,
    24'b100100010010000000100101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000110000101011,
    24'b000001100011000101100001,
    24'b001000110101111110101100,
    24'b000010100110011111000011,
    24'b000001010110100011001111,
    24'b000000010110011011010101,
    24'b000000010110100011001111,
    24'b000000000110011011010011,
    24'b000000000110011111001111,
    24'b000000000110011111001100,
    24'b000000000110011111001101,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011011010011,
    24'b000000000110011111001110,
    24'b000000000110011011010010,
    24'b000000000110011011010100,
    24'b000000010110010111010011,
    24'b000000000110011111010001,
    24'b000000000110100011010000,
    24'b000000000110010111001100,
    24'b000010000110010111001101,
    24'b000000100110010111010001,
    24'b000010000110011011001100,
    24'b000111000110001010111000,
    24'b000110100011111001111111,
    24'b000000010001010100111101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010100110000001100000011,
    24'b101011000010000100101000,
    24'b110011100010100100101111,
    24'b111000010010000000100111,
    24'b111011100001101000100110,
    24'b111010100001110000100100,
    24'b111010110001110000100100,
    24'b111011000001101100100100,
    24'b111011010001101100100100,
    24'b111011000001101000100100,
    24'b111011010001101100100100,
    24'b111011010001101100100100,
    24'b111010100001110100100011,
    24'b111011100001101100100101,
    24'b110111010010001100101010,
    24'b110010000010100000101110,
    24'b101001010010000000101001,
    24'b001100100000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000101100101101,
    24'b000001100010010101011101,
    24'b000110000101110010100101,
    24'b000010010110000110111100,
    24'b000010000110100111001111,
    24'b000001000110010111001110,
    24'b000001010110011011001100,
    24'b000000010110011111001101,
    24'b000000000110011111001101,
    24'b000000000110011011010011,
    24'b000000010110011011010000,
    24'b000000010110011011001110,
    24'b000000000110011111001111,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000100110100111010010,
    24'b000000000110011111010000,
    24'b000000010110011011001101,
    24'b000000010110011011010010,
    24'b000000100110011011010010,
    24'b000001000110010111001110,
    24'b000010000110011011001000,
    24'b000010110110001111000001,
    24'b000111110110011110111010,
    24'b000110010100101110001011,
    24'b000001010010000001001011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001011010000000000000001,
    24'b010001100000011000000010,
    24'b101100100010111100110110,
    24'b101011000011000000110101,
    24'b101011000011000000110101,
    24'b101011000011000000110101,
    24'b101010110011000000110100,
    24'b101011000011000000110101,
    24'b001101100000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001011000111001,
    24'b000011010011100001101111,
    24'b000111000101100110100101,
    24'b000101000110010011000001,
    24'b000001000110000011000011,
    24'b000000100110001111001010,
    24'b000001000110100011001111,
    24'b000001100110100011010100,
    24'b000000110110011111010110,
    24'b000000010110011111010010,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011011001101,
    24'b000000000110011011010010,
    24'b000000000110011011010100,
    24'b000000010110011011010010,
    24'b000000110110011011001110,
    24'b000000010110110111010000,
    24'b000000110110110011001111,
    24'b000011100110011111001001,
    24'b000110010110000110111010,
    24'b001000100101111010101001,
    24'b000011100100010110000100,
    24'b000010100010101101011000,
    24'b000000000001000100110011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001000100110010,
    24'b000000000001111101001010,
    24'b000010000011010001101001,
    24'b000101000101001110010101,
    24'b000101100110001110111101,
    24'b000100100110011111000101,
    24'b000010100110100011001010,
    24'b000000000110001111001001,
    24'b000000000110011111001110,
    24'b000000010110011111001101,
    24'b000000110110011011001110,
    24'b000000110110011011010010,
    24'b000000110110100011010100,
    24'b000000010110011111010010,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010011,
    24'b000000000110011011010100,
    24'b000000000110011011010011,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000010110100111001110,
    24'b000000100110100011001101,
    24'b000001000110010111001101,
    24'b000001100110010011010000,
    24'b000010000110010011000111,
    24'b000011110110000110111001,
    24'b000101000101111010100111,
    24'b000110000101011010010111,
    24'b000011010100100110000011,
    24'b000100110011110101111010,
    24'b000100000011100101110101,
    24'b000011010011100001101110,
    24'b000011110011101101101111,
    24'b000011100011110001110010,
    24'b000101000100010001111111,
    24'b000101110101000110011000,
    24'b000110100101100110100110,
    24'b000101100101110110110000,
    24'b000100000110000110111001,
    24'b000010010110010011000010,
    24'b000001110110010111001011,
    24'b000001000110010111001111,
    24'b000000100110010111001101,
    24'b000000010110011011001101,
    24'b000000110110011011001100,
    24'b000000100110011011001100,
    24'b000000110110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011010001,
    24'b000000010110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010100,
    24'b000000100110010111010001,
    24'b000000100110010111010000,
    24'b000000010110011011010001,
    24'b000000010110011111010001,
    24'b000000000110011111001110,
    24'b000000000110011011001101,
    24'b000001000110011011000110,
    24'b000000110110010111000111,
    24'b000001010110010011001001,
    24'b000000100110011111001000,
    24'b000010000110100011000110,
    24'b000010100110100011000101,
    24'b000010100110011011000100,
    24'b000010010110011011000001,
    24'b000010010110010110111111,
    24'b000010000110011111000010,
    24'b000001100110010111000011,
    24'b000001000110010011000110,
    24'b000001010110011011001011,
    24'b000000110110100011001100,
    24'b000000110110100011001010,
    24'b000000100110011111001100,
    24'b000000100110011011001111,
    24'b000000010110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010010,
    24'b000000100110011011010010,
    24'b000000010110011011001111,
    24'b000000010110011011001110,
    24'b000000000110011011010001,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001111,
    24'b000000010110011011001111,
    24'b000000010110011011001111,
    24'b000000010110011111001111,
    24'b000000010110011011010001,
    24'b000000010110011111010000,
    24'b000000100110011011010001,
    24'b000000010110011011010011,
    24'b000000000110011011010010,
    24'b000000000110011111001111,
    24'b000000010110100011001111,
    24'b000000000110100011001111,
    24'b000000010110011111010000,
    24'b000000000110011011001111,
    24'b000000010110011111001111,
    24'b000000100110011011010001,
    24'b000000110110011011010010,
    24'b000001000110011111001110,
    24'b000001010110011111001110,
    24'b000001010110011011001110,
    24'b000000110110010111001100,
    24'b000000110110011011001101,
    24'b000000110110011011001111,
    24'b000000100110011111010010,
    24'b000000010110100011010101,
    24'b000000010110011111010010,
    24'b000000000110011111010000,
    24'b000000100110011011010010,
    24'b000000010110011111001111,
    24'b000000010110011011010010,
    24'b000000000110011011010011,
    24'b000000010110011011010011,
    24'b000000010110011011001111,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000100110011111010100,
    24'b000000000110011011010011,
    24'b000000110110010111010010,
    24'b000000110110010111010000,
    24'b000001000110011011010001,
    24'b000000110110010111010010,
    24'b000000100110011011010011,
    24'b000000010110011011010010,
    24'b000000010110011011001111,
    24'b000000010110011011001101,
    24'b000000000110011111001011,
    24'b000000000110011111001110,
    24'b000000010110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011011010001,
    24'b000000000110011111010010,
    24'b000000010110011111010011,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011011010000,
    24'b000000100110010111010000,
    24'b000000010110011011010010,
    24'b000000010110011111010101,
    24'b000000010110011011010010,
    24'b000000010110011011001111,
    24'b000000010110011111001011,
    24'b000000000110100011001011,
    24'b000000000110011111001111,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000010110100111001111,
    24'b000000100110100111010010,
    24'b000000100110100111010010,
    24'b000000010110011111010011,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000100110100011010100,
    24'b000000000110100111010110,
    24'b000000100110011111010011,
    24'b000000010110011011010000,
    24'b000000010110100011001101,
    24'b000000010110100011001101,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000
};


assign mem_red = memory_red;

logic [23:0] memory_green [0:4899] = '{
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011001111,
    24'b000000010110100011001111,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010011,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000010110100011010001,
    24'b000000000110010111010001,
    24'b000000010110011011010010,
    24'b000000010110010111010011,
    24'b000000010110010111010011,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011001111,
    24'b000000000110011011001111,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000010110011111010010,
    24'b000000000110011011010001,
    24'b000000000110011111001111,
    24'b000000100110011011001110,
    24'b000000100110011011001110,
    24'b000000100110010111010000,
    24'b000000100110011011001110,
    24'b000000100110011011001110,
    24'b000000000110011111001101,
    24'b000000010110100011001101,
    24'b000000000110011111001100,
    24'b000000010110100011001101,
    24'b000000000110011111001110,
    24'b000000000110011111001101,
    24'b000000000110011111001100,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011001111,
    24'b000000010110100011001111,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110100011010011,
    24'b000000000110100011010011,
    24'b000000000110100011010011,
    24'b000000000110100011010011,
    24'b000000000110011111010011,
    24'b000000000110011011010010,
    24'b000000010110011011010001,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000010110100011010000,
    24'b000000100110100111010001,
    24'b000000010110100011001111,
    24'b000000000110011111001111,
    24'b000000000110011111001101,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000100110011111001110,
    24'b000000010110011011001111,
    24'b000000100110011111010011,
    24'b000000100110011011010100,
    24'b000000100110011011010101,
    24'b000000000110100011010010,
    24'b000000000110100011010010,
    24'b000000000110100011010000,
    24'b000000010110100011001111,
    24'b000000100110100011001111,
    24'b000000100110100011010000,
    24'b000000100110011011010001,
    24'b000000010110011111001110,
    24'b000000010110011011001101,
    24'b000000110110100011010001,
    24'b000001000110100011010100,
    24'b000001010110100111010100,
    24'b000000110110011111010010,
    24'b000000110110011111010010,
    24'b000000100110011011010011,
    24'b000000100110011111010100,
    24'b000000100110011111010100,
    24'b000000100110011111010001,
    24'b000000100110011111010010,
    24'b000000100110011111010010,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001101,
    24'b000000000110011011001011,
    24'b000000000110010111001110,
    24'b000000010110011011010010,
    24'b000000010110010111010100,
    24'b000000000110010011010100,
    24'b000000010110100011001110,
    24'b000000100110011111001100,
    24'b000001010110011111001100,
    24'b000001100110010111001001,
    24'b000010000110010011000111,
    24'b000010000110010011000110,
    24'b000010010110010111001000,
    24'b000001110110010011000010,
    24'b000010000110011011000010,
    24'b000010000110010111000100,
    24'b000010010110010111001000,
    24'b000001010110010011000111,
    24'b000001010110011011001000,
    24'b000001010110010111001011,
    24'b000001010110011011001110,
    24'b000000110110010111001111,
    24'b000000110110010111010001,
    24'b000000100110011111010001,
    24'b000000100110011111010001,
    24'b000001000110011011010001,
    24'b000000100110011111010001,
    24'b000000000110010111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100011010001,
    24'b000000000110011111010000,
    24'b000000100110011011010001,
    24'b000000010110100011010001,
    24'b000000010110011011001111,
    24'b000000000110010111001111,
    24'b000000010110011011010000,
    24'b000001100110101111010101,
    24'b000001100110011111010101,
    24'b000000110110010111001101,
    24'b000001100110010111001000,
    24'b000011000110010011000011,
    24'b000011110110001010111101,
    24'b000101000110001110111011,
    24'b000101100110000110110110,
    24'b000101100101110010101111,
    24'b000101010101100110101011,
    24'b000101000101101110100110,
    24'b000100110101101110100101,
    24'b000100100101101110100111,
    24'b000101110101111010110000,
    24'b000101000110001110110111,
    24'b000011000110000010111000,
    24'b000010100110010010111101,
    24'b000010100110010111000010,
    24'b000001100110001111000110,
    24'b000001110110010111001110,
    24'b000001100110011011001101,
    24'b000000100110100111001101,
    24'b000001100110100011010001,
    24'b000000110110010111010001,
    24'b000000010110100011001111,
    24'b000000000110011111010011,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110100011010000,
    24'b000000000110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010000,
    24'b000000010110011111010101,
    24'b000000110110010111001111,
    24'b000000000110011011001010,
    24'b000000000110011111001101,
    24'b000001000110100111010011,
    24'b000000110110001111001011,
    24'b000100000110100011000111,
    24'b000010110110001010111010,
    24'b000101000110011011000001,
    24'b000110110110000110110001,
    24'b001000010101101110011110,
    24'b000100010100000001111010,
    24'b000010010010011101010110,
    24'b000000000001100100111101,
    24'b000000000001000100101100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001011000110101,
    24'b000000000001111001001010,
    24'b000010100010111101101001,
    24'b000111000101010010010001,
    24'b000110110101110110100110,
    24'b000101110101111010110100,
    24'b000011110110010011000010,
    24'b000010000110010011001110,
    24'b000001100110011111001100,
    24'b000000100110110011001111,
    24'b000001010110010011010000,
    24'b000000110110010011010101,
    24'b000000000110011111010001,
    24'b000000000110100011001100,
    24'b000000100110011111001111,
    24'b000000100110011011010001,
    24'b000000010110011011001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000110110010111010000,
    24'b000000010110011011001101,
    24'b000000010110100111001011,
    24'b000001100110011011001101,
    24'b000011000110010111001000,
    24'b000100110110001110111110,
    24'b001000000101111110101100,
    24'b000111110100110110001100,
    24'b000001110010001101011000,
    24'b000000010001001000110011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001111011001000001010111,
    24'b010000001001001101010000,
    24'b001000101010110101001110,
    24'b001000011011000001001011,
    24'b001000111011001001001011,
    24'b001001111011001001001100,
    24'b001001101010111101001100,
    24'b001001101010110001001100,
    24'b001101101001101001010110,
    24'b010000101000111101011110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000100001010100110111,
    24'b000100010011100001110101,
    24'b001001010101100010101001,
    24'b000101100110100111000110,
    24'b000010110110010011000101,
    24'b000010000110011011001000,
    24'b000001000110010011001101,
    24'b000001010110011111001100,
    24'b000000100110011011001010,
    24'b000000100110010011001110,
    24'b000000100110010111010010,
    24'b000000000110011011010011,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000001000110011011001110,
    24'b000001000110100011001101,
    24'b000000110110010011010101,
    24'b000000110110011111011000,
    24'b000010000110001011000010,
    24'b000111100101101110101111,
    24'b000010110011101001111011,
    24'b000000010001010000111110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001011101000001001000111,
    24'b001011111010100001010101,
    24'b001000101011000001010000,
    24'b001000101011000101001110,
    24'b001001011010111101001111,
    24'b001000101011000101001110,
    24'b001000111011000001001101,
    24'b001000111011000101001111,
    24'b001000101011000101001111,
    24'b001001001011000001001111,
    24'b001001001011000001001111,
    24'b001001001011000001001111,
    24'b001001101010111101001100,
    24'b001000101011000001001110,
    24'b001001001011000001010000,
    24'b001001011010111001010010,
    24'b001101001010011001010110,
    24'b001011011000010001000111,
    24'b000000000000000000000000,
    24'b000000010000111100101000,
    24'b000010000010001001010110,
    24'b000111100100100010010100,
    24'b000100100110001110110110,
    24'b000010010110100111001000,
    24'b000000110110011011001010,
    24'b000000010110001111001101,
    24'b000000010110011111010101,
    24'b000001000110101111011001,
    24'b000000100110001111010010,
    24'b000000010110011011010000,
    24'b000000100110011111010001,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010000,
    24'b000000000110011111010000,
    24'b000000100110011111001011,
    24'b000001110110100011000110,
    24'b000011010110011011000111,
    24'b000100100101110110110110,
    24'b000011110011110001111001,
    24'b000001000001000000110100,
    24'b000000000000000000000000,
    24'b001011000111000000111011,
    24'b001011101010110101010010,
    24'b001001111011000001001011,
    24'b001001001011000101010000,
    24'b001000101011000101001101,
    24'b001001001011000001001011,
    24'b001000111011000101001010,
    24'b001000101011000101001110,
    24'b001001001011000001001100,
    24'b000111011011010001001011,
    24'b001001001011000001001101,
    24'b001000111011000101001101,
    24'b001000101011000101001101,
    24'b001000011011001001001101,
    24'b001000001011001101001011,
    24'b000111101011001101001110,
    24'b001000011011000101001100,
    24'b001001001011000101001001,
    24'b001000011011001001001010,
    24'b001000011011000101001110,
    24'b001000101011000001010001,
    24'b001010001010111001010101,
    24'b001010011010101001010011,
    24'b001000100101100000110001,
    24'b000000000000000000000000,
    24'b000001110010010001010001,
    24'b000101010101011110100000,
    24'b000100000110011110111110,
    24'b000010000110110011010001,
    24'b000001010110010011010001,
    24'b000010010110000111001011,
    24'b000001110110010011001010,
    24'b000000110110011011001110,
    24'b000000110110010111010000,
    24'b000000010110011011010000,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000010110100011010001,
    24'b000000010110011111010001,
    24'b000001010110011011001100,
    24'b000101100110001110111111,
    24'b000110000100111010010010,
    24'b000000100001010100111001,
    24'b000000000000000000000000,
    24'b000110110110000000110000,
    24'b001100001010101101010010,
    24'b001000111011010001001101,
    24'b001000101011000101001111,
    24'b001000011011000001001001,
    24'b001000111011000001001101,
    24'b001000111011000001001111,
    24'b001000111011000101001011,
    24'b001001101010111101001100,
    24'b000111111011001101001110,
    24'b001001011011000001001101,
    24'b001000111011001001001010,
    24'b001000111011000101001100,
    24'b001000111011000101001110,
    24'b001000111011000101001110,
    24'b001001001011000101001101,
    24'b001001001011001001001010,
    24'b001000111011000101001101,
    24'b001000101011000101001101,
    24'b001000111011000101001110,
    24'b001000101011001001010000,
    24'b001000111011000001001110,
    24'b001000101011001001001011,
    24'b001000101011001001001110,
    24'b001001011010111101001110,
    24'b001001001011001001001001,
    24'b001100101010011101011000,
    24'b001000110101011100111000,
    24'b000000000000000000000000,
    24'b000011100011010001100100,
    24'b000110110110000110110000,
    24'b000011110110010111001010,
    24'b000001110110010011001110,
    24'b000000110110100011010001,
    24'b000000110110011011001110,
    24'b000000100110010111001101,
    24'b000000010110011011010000,
    24'b000000100110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011010000,
    24'b000000000110011011010011,
    24'b000000100110011111010000,
    24'b000000010110011011001101,
    24'b000000000110100011010011,
    24'b000001010110011011010111,
    24'b000001000110011111010000,
    24'b000011100110011011000101,
    24'b000110010110000110110001,
    24'b000011010011011001110000,
    24'b000000000000000000000000,
    24'b000110110100001000100010,
    24'b001100011010100101010110,
    24'b001001001010111101010000,
    24'b001000111011000101001100,
    24'b001000111011000101001100,
    24'b001000011011000101001110,
    24'b001000111011000101001101,
    24'b001000111011000001001101,
    24'b001000101011000101001101,
    24'b001000101011000101001101,
    24'b001000111011000001001101,
    24'b001000011011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000001001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000011011000101001110,
    24'b001000111011000101001101,
    24'b001000111011000101001011,
    24'b001000111011000101001101,
    24'b001000111011000001001101,
    24'b001000111011000101001100,
    24'b001000011011000101001101,
    24'b001001011010111101001111,
    24'b001110001010010101011001,
    24'b000000000000000000000000,
    24'b000000100001100101000001,
    24'b001000000101011010100010,
    24'b000011100110011011000100,
    24'b000001110110100111001111,
    24'b000001000110101011010100,
    24'b000000010110011011010001,
    24'b000001000110010111010001,
    24'b000001010110011111010010,
    24'b000000100110010111001101,
    24'b000000010110011011001110,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011010000,
    24'b000000000110011011010011,
    24'b000000010110011011010000,
    24'b000000000110100111001101,
    24'b000000010110011011001101,
    24'b000000010110100011001110,
    24'b000001100110011011000001,
    24'b000110010101110010101011,
    24'b000001010010010001010100,
    24'b000000000000000000000000,
    24'b000101100101010100100011,
    24'b001010001011001101010001,
    24'b001000111010111101001001,
    24'b001000101011000001001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001001011011001001010001,
    24'b001011101010111001010011,
    24'b000011010011001000010111,
    24'b000000000001010000101011,
    24'b000101100100010101111110,
    24'b000111000110011110111110,
    24'b000001100110011111001110,
    24'b000010010110001111001011,
    24'b000000100110011111001100,
    24'b000001000110100011010001,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000100110011111010001,
    24'b000001100110001111010000,
    24'b000000000110100011010000,
    24'b000001010110010111001100,
    24'b000011010101110110111001,
    24'b000101110101011010010110,
    24'b000001000001010101000101,
    24'b000000000000000000000000,
    24'b001111001010000101011100,
    24'b000111111011000101001110,
    24'b001000111011001101001100,
    24'b001001011011010101001100,
    24'b001001011011000001001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001001001011001001010000,
    24'b001000001011000001000101,
    24'b000111111011000001001010,
    24'b001010110111001100111110,
    24'b000000000000000000000000,
    24'b000100010011101001110100,
    24'b000011010110011010111000,
    24'b000011110110000111001000,
    24'b000000100110001111010000,
    24'b000000110110100111010011,
    24'b000000000110100111001110,
    24'b000000110110010111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010011,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110010111001111,
    24'b000000010110010111010000,
    24'b000000100110011111010001,
    24'b000000000110100011010001,
    24'b000001010110011011010000,
    24'b000011110110001111000101,
    24'b001000110110000010100101,
    24'b000000000000110000101011,
    24'b000000000000000000000000,
    24'b001110111001110101010101,
    24'b000110101011010101001011,
    24'b001010001010110101001111,
    24'b001001001010111101010010,
    24'b001000001011001001001101,
    24'b001000101011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111010111101010011,
    24'b001001001011000101001011,
    24'b001001001010111101001111,
    24'b001001101011000001010000,
    24'b001101101010001101010110,
    24'b000000000000000000000000,
    24'b000100110011100001101100,
    24'b000110000110010110111110,
    24'b000001010110011111010110,
    24'b000001010110101011010010,
    24'b000000110110011011001101,
    24'b000000010110011011010001,
    24'b000000000110011111001110,
    24'b000000010110100011001111,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110010111010001,
    24'b000000110110100011010010,
    24'b000001000110011111001110,
    24'b000000100110100011001011,
    24'b000010000110010111000010,
    24'b000111010101111110100101,
    24'b000000000001010100110101,
    24'b000000000000000000000000,
    24'b001100011010100001010110,
    24'b001010001010110101001101,
    24'b001001011011001001001000,
    24'b001000001011001001001010,
    24'b001000011011001001001010,
    24'b000111111011001001001101,
    24'b001000111011000001001111,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001001001011000001001100,
    24'b000111111011001001001111,
    24'b001001111010111001001111,
    24'b001000111011000001000111,
    24'b001000101011001001001100,
    24'b001110011010010101010111,
    24'b000000000000000000000000,
    24'b000011010011110101101110,
    24'b000100000110011110111101,
    24'b000010100110010111001010,
    24'b000001010110010111001111,
    24'b000000000110100011010011,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010011,
    24'b000000100110011011001111,
    24'b000001010110011111001110,
    24'b000001100110011011000111,
    24'b000111010110000010101110,
    24'b000000100001001101000000,
    24'b000000000000000000000000,
    24'b001101001001100101010001,
    24'b001000011011000101001110,
    24'b000111111011001001001011,
    24'b001000001011000101001101,
    24'b001001001010111101010001,
    24'b001000011011001001001010,
    24'b001001001011000001001011,
    24'b001000111011000101001110,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000011011001001001101,
    24'b001000101011000101001011,
    24'b001000001011001101001011,
    24'b001000111011000001010010,
    24'b001001001011000101010000,
    24'b001000011011000101001000,
    24'b001011010111011100111111,
    24'b000000000000000000000000,
    24'b000110000100111010000110,
    24'b000101010101111110111110,
    24'b000001010110010011010001,
    24'b000000010110011011010100,
    24'b000000010110011111010101,
    24'b000000000110011011010010,
    24'b000000000110011111010001,
    24'b000000000110011111001110,
    24'b000000000110011111001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010010,
    24'b000000010110011011001111,
    24'b000000100110011011001101,
    24'b000000000110100011010100,
    24'b000001110110100111010000,
    24'b000010000110001111000111,
    24'b000101010110010010111100,
    24'b000010010010101001011101,
    24'b000000000000000000000000,
    24'b001111111001101101011000,
    24'b001000101011001001001001,
    24'b001000111011000101010000,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001010001010111001001111,
    24'b001001110110100100111000,
    24'b000000000001010000101101,
    24'b000111110101100110011111,
    24'b000100110110100011000101,
    24'b000000110110011111010011,
    24'b000001010110100011010101,
    24'b000000010110010111010101,
    24'b000000010110011011010010,
    24'b000000010110011111001110,
    24'b000000010110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001100,
    24'b000000000110100011001011,
    24'b000000010110100011010000,
    24'b000000010110001111001010,
    24'b000011100110000110110110,
    24'b000100010100000101110111,
    24'b000000000000000000000000,
    24'b000110100101001100100011,
    24'b000111011011001001001101,
    24'b001000011010111101001011,
    24'b001000101011000001001010,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000011011000001001100,
    24'b001010101010111001001110,
    24'b000000000000000000000000,
    24'b000001000001101001000000,
    24'b000110110110000010101111,
    24'b000010100110011011001001,
    24'b000000100110001111010001,
    24'b000001000110011011010001,
    24'b000000110110010111010000,
    24'b000000100110010111010010,
    24'b000000010110011111010101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010000,
    24'b000000010110011111010011,
    24'b000000010110011111010000,
    24'b000001010110011011010010,
    24'b000010100110010011001010,
    24'b000110100101101010100000,
    24'b000000000001001100101101,
    24'b000000000000000000000000,
    24'b001001111010110101001111,
    24'b001001001010111001001100,
    24'b001000101011001001001101,
    24'b001000101011000001001011,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000101011000001001100,
    24'b001001101011000001001010,
    24'b001011001010101101010010,
    24'b000000000000000000000000,
    24'b000010100011001101101101,
    24'b000010100110000010111011,
    24'b000001110110100011010101,
    24'b000000000110011111001111,
    24'b000000110110011011001110,
    24'b000001000110010111001111,
    24'b000000010110011111010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110010111010100,
    24'b000000110110010011010101,
    24'b000001100110001011010000,
    24'b000110000110000110111010,
    24'b000001110010101001011100,
    24'b000000000000000000000000,
    24'b001110111010001101010111,
    24'b001000101011001101010000,
    24'b001000111011000001010000,
    24'b000111111011001101001001,
    24'b001001001011000001001111,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000011011000101001111,
    24'b001001001010111101001111,
    24'b001001001011000001001101,
    24'b000111110110001000101110,
    24'b000000000000000000000000,
    24'b001000000101110110100100,
    24'b000010100110011111000110,
    24'b000000000110011011010010,
    24'b000000100110011111010001,
    24'b000001000110011011001011,
    24'b000000010110011011001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000110110011011001100,
    24'b000001010110010011010010,
    24'b000010010110001111001001,
    24'b000111010101010110010101,
    24'b000000000000000000000000,
    24'b000110000101000100100010,
    24'b001001011011000001001110,
    24'b001001001011000101001011,
    24'b000111101011001101001101,
    24'b001000101011000101001011,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000011011000101001111,
    24'b000111111011001001001101,
    24'b000111111011001001001111,
    24'b001000101011001001001111,
    24'b000000000000000000000000,
    24'b000001010010100001001110,
    24'b000110110110011010110100,
    24'b000001110110011011010011,
    24'b000000100110011111010100,
    24'b000001000110100011001010,
    24'b000000000110011111010010,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000010110011111001111,
    24'b000000100110011111010011,
    24'b000000010110011011010010,
    24'b000000110110100011001100,
    24'b000000110110000111001011,
    24'b000101000110001110111101,
    24'b000001100010011001001100,
    24'b000000000000000000000000,
    24'b001010111010101101010010,
    24'b001000101011000101001100,
    24'b001000101011000101001100,
    24'b001001001011000001001100,
    24'b001000111011000001001101,
    24'b001000101011000101001100,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001001011010111101001111,
    24'b001000111011000101001010,
    24'b001000011011001001001111,
    24'b001001011010111101001100,
    24'b001011101001101101010100,
    24'b000000000000000000000000,
    24'b001001100110000010100000,
    24'b000001010101110011000110,
    24'b000001100110011011001110,
    24'b000001000110100011010011,
    24'b000000000110100011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000010110011111001101,
    24'b000001000110011011010011,
    24'b000000110110010111010011,
    24'b000001000110011011001000,
    24'b000100110110110011010000,
    24'b000111100101110110100100,
    24'b000000000000000000000000,
    24'b001000100101011100101111,
    24'b001001011010111101001110,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001110,
    24'b001000111011000101001011,
    24'b000111111011001001001110,
    24'b001001101011000101001011,
    24'b001001111010111001010010,
    24'b000000000000000000000000,
    24'b000000110010001001010100,
    24'b000101010110011111000011,
    24'b000010010110010111001001,
    24'b000000000110011111010011,
    24'b000000000110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111001111,
    24'b000000110110010111010010,
    24'b000000110110010111010001,
    24'b000001000110100011000101,
    24'b000100100101111110110101,
    24'b000001110010101101011010,
    24'b000000000000000000000000,
    24'b001110111010001101010010,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000001001110,
    24'b001000101011000101001110,
    24'b001000111011000001000111,
    24'b001001001011000001001001,
    24'b001011001000011101001000,
    24'b000000000000000000000000,
    24'b001000000110000010101010,
    24'b000011000110010011001011,
    24'b000000000110011111010001,
    24'b000000100110010111001100,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000110110010111010010,
    24'b000000110110010111010000,
    24'b000000100110100011001001,
    24'b000110000110100010110000,
    24'b000000000000101100101100,
    24'b000000000000000000000000,
    24'b001000011011000101001100,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001010,
    24'b001000111011000101001111,
    24'b001000111011000101001111,
    24'b001000011011001001001101,
    24'b001000011011001001001100,
    24'b001100001010100001010010,
    24'b000000000000000000000000,
    24'b000111110100010101111111,
    24'b000011110110001011000110,
    24'b000000000110011011010010,
    24'b000000110110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110010111010100,
    24'b000000110110010111010001,
    24'b000000010110011111001110,
    24'b000001110110011111001000,
    24'b000111110101010110010110,
    24'b000000000000000000000000,
    24'b001011100111000000111011,
    24'b001000001011000001001010,
    24'b001000011011001001001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011001001001001,
    24'b001000101011000101001111,
    24'b001000111011000101001100,
    24'b001000101011000101001111,
    24'b001000011011001001010000,
    24'b001010011010111001001101,
    24'b000100010011000100010100,
    24'b000000000001010100111110,
    24'b000110100110010010111011,
    24'b000001010110011011001111,
    24'b000000010110011111010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011011010001,
    24'b000000000110010111010101,
    24'b000000110110010111010000,
    24'b000000110110011111001000,
    24'b000100010110010111000100,
    24'b000001100010101001100001,
    24'b000000000000000000000000,
    24'b001100011010100101001110,
    24'b001000101011000001001010,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000011011001001001101,
    24'b001000101011000101001111,
    24'b001000111011001001001000,
    24'b001001101010111101001101,
    24'b001000101011000101001111,
    24'b001000011011001001000111,
    24'b010000011000111101010110,
    24'b000000000001010000101100,
    24'b000111000110000110100111,
    24'b000001100110010111001010,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010001,
    24'b000000110110011011001110,
    24'b000000110110011011001100,
    24'b000011110110001010111000,
    24'b000000010001001100110011,
    24'b000000000000000000000000,
    24'b001010101010110101001010,
    24'b001000011011000001001101,
    24'b001000111011000101001110,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001100,
    24'b001001001011000101010001,
    24'b000000000000000000000000,
    24'b000111010101011010010000,
    24'b000010110110010111001010,
    24'b000000110110011111010001,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010000,
    24'b000000110110010111001111,
    24'b000001010110010111001011,
    24'b000101010101110010101001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001001111011000001001010,
    24'b001001001011000101001011,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000101011000001001100,
    24'b001000111011000001001110,
    24'b000000000000000000000000,
    24'b000011100011110101110000,
    24'b000011110110010111000100,
    24'b000000010110011011001111,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010000,
    24'b000000110110010111010000,
    24'b000010000110010011001011,
    24'b001000110101111010100010,
    24'b000000000000000000000000,
    24'b001100001000001001000111,
    24'b001000111011000101001100,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001001011011000101001100,
    24'b000000000000000000000000,
    24'b000000100001111101001001,
    24'b000100110110001110111001,
    24'b000000100110011011001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001111,
    24'b000000110110010111010000,
    24'b000010010110001111001010,
    24'b001000100101001010001110,
    24'b000000000000000000000000,
    24'b001011011000010101000100,
    24'b001000011011000101001111,
    24'b001000111011000101010000,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000101011000101001100,
    24'b001000001011000001001010,
    24'b000001000010100100000110,
    24'b000000000001001100110101,
    24'b000101000110000110110010,
    24'b000000110110011011001110,
    24'b000000010110011011010001,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011011001111,
    24'b000000100110010111010000,
    24'b000010100110010111001001,
    24'b000110100100001101110110,
    24'b000000000000000000000000,
    24'b001110101010001101010110,
    24'b001000101011000101001100,
    24'b001000101011000101001111,
    24'b001000111011000001001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001001011011001001001100,
    24'b001110011010000101011110,
    24'b000000000000101100101101,
    24'b000101110110000110110001,
    24'b000001000110011011001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111001111,
    24'b000000010110011111001111,
    24'b000000110110010111001111,
    24'b000011000110010111000110,
    24'b000011010011010001100010,
    24'b000000000000000000000000,
    24'b001100101010100001010100,
    24'b001000101011001001001010,
    24'b001001001011000001001011,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000101011001101001110,
    24'b001110001010001101011001,
    24'b000000000000101000101011,
    24'b000110100110000110101111,
    24'b000001000110010111001110,
    24'b000000010110011011010001,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111001110,
    24'b000001100110011111010000,
    24'b000011110110010111000111,
    24'b000001110010110101011110,
    24'b000000000000000000000000,
    24'b001101011010011001010100,
    24'b001001001011000101001100,
    24'b001000111011000101001010,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000011011001001001101,
    24'b001110101010001001010100,
    24'b000000000000000000000000,
    24'b000110100101111110101011,
    24'b000001000110011011001111,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010000,
    24'b000001100110011111010010,
    24'b000011000110011011001001,
    24'b000001110010100101011101,
    24'b000000000000000000000000,
    24'b001101011010011101010010,
    24'b001001011011000001001101,
    24'b001000111011000001001110,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001001001011000001001101,
    24'b001000001011001001001101,
    24'b001111001010000101010110,
    24'b000000000000000000000000,
    24'b000101100110000110101101,
    24'b000000100110011011001110,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000010110011111010001,
    24'b000001100110011111010010,
    24'b000011100110010111001001,
    24'b000010100010110101100001,
    24'b000000000000000000000000,
    24'b001100011010100001010001,
    24'b001000001011001001001101,
    24'b001001001011000001001110,
    24'b001000111011000101001110,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000001001101,
    24'b001000011011000001001011,
    24'b001101001010010001010111,
    24'b000000010000011100101010,
    24'b000110000101111110101101,
    24'b000001000110011011001110,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010001,
    24'b000001010110011011010010,
    24'b000011100110010111001001,
    24'b000011110011110001101111,
    24'b000000000000000000000000,
    24'b001101101010010101010101,
    24'b000111011011001101001110,
    24'b001001001011000001001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000101011000101001101,
    24'b001000111011000101001111,
    24'b001111011010000001011100,
    24'b000000000000101100110001,
    24'b000110100101111010110000,
    24'b000001010110011011010000,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010011,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000100110011111001111,
    24'b000001100110011111001111,
    24'b000010100110010011000101,
    24'b000111000101001010000011,
    24'b000000000000000000000000,
    24'b001011001000010101000101,
    24'b001001001011000001001111,
    24'b001000011011001101001010,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000101011000101001100,
    24'b001000011011000101010000,
    24'b000001010010100100000110,
    24'b000000000001000100111000,
    24'b000100110110001110110100,
    24'b000000100110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111001111,
    24'b000000010110011111001100,
    24'b000001000110010011000100,
    24'b000111100101100010010101,
    24'b000000000000000000000000,
    24'b001100001000001101000100,
    24'b001000011011000001001110,
    24'b001000101011001001001010,
    24'b001000101011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000011011001001001010,
    24'b001000101010111001001110,
    24'b000000000000000000000000,
    24'b000000000001011001000001,
    24'b000011000110001110111000,
    24'b000000000110100111001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011111001111,
    24'b000000100110011111001101,
    24'b000001000110010011001000,
    24'b000111010101111110100110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001001101011000001001110,
    24'b001000111011000001001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001001001010111101001111,
    24'b000000000000000000000000,
    24'b000010100011001101100001,
    24'b000011010110001010111111,
    24'b000001110110010011001111,
    24'b000000100110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000100110011111001111,
    24'b000000110110010111001100,
    24'b000101100110000010110010,
    24'b000000000001000100110000,
    24'b000000000000000000000000,
    24'b001001101010111101001010,
    24'b001001001010111101001111,
    24'b001000111011000101001110,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001001111010111101001111,
    24'b000000000000000000000000,
    24'b001000010100110110000110,
    24'b000011000110000111000110,
    24'b000000010110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011001111,
    24'b000000000110011111001110,
    24'b000000100110011111001111,
    24'b000000000110010011001100,
    24'b000101010110000110111001,
    24'b000000100010000101001000,
    24'b000000000000000000000000,
    24'b001100011010111101010010,
    24'b001000101011000101001100,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001001001011001001001110,
    24'b010000001001010001010001,
    24'b000000000000000000000000,
    24'b001000010101100010011111,
    24'b000010110110010111001011,
    24'b000000010110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111001110,
    24'b000000010110100011001101,
    24'b000000000110011011001101,
    24'b000000010110010111001111,
    24'b000000110110100111010010,
    24'b000100000110010111000011,
    24'b000101110100101110000011,
    24'b000000000000000000000000,
    24'b001011010110111000111010,
    24'b001000101011000001001100,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001001001010111101001111,
    24'b000011110011001100010110,
    24'b000000000000100100110011,
    24'b001000110110000010111100,
    24'b000001010110100111001010,
    24'b000000100110010011001111,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111001110,
    24'b000000000110011111001100,
    24'b000000000110011011001101,
    24'b000000000110010011001110,
    24'b000001100110101011010100,
    24'b000001100110011011001000,
    24'b000111110110001110101001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001001101010111001001110,
    24'b001000111011000101001101,
    24'b001000111011000001001101,
    24'b001000111011000101001011,
    24'b001000011011000101001101,
    24'b001000111011000101001110,
    24'b001000111011000101001011,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000011011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001100,
    24'b001000111011000001001101,
    24'b001101101010011001010000,
    24'b000000000000000000000000,
    24'b000011110010101101011110,
    24'b000100000110001111000110,
    24'b000001000110101011010001,
    24'b000000010110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000001010110100111010010,
    24'b000000100110100011010000,
    24'b000101100110100010111110,
    24'b000001010001110001001110,
    24'b000000000000000000000000,
    24'b001101111010011001010100,
    24'b001001001011000101001100,
    24'b001000101011000101001110,
    24'b001000111011001001001000,
    24'b001000101011001001001101,
    24'b001001001010111101010010,
    24'b001000101011001001001000,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000001011001001001100,
    24'b001001001011000001001101,
    24'b001000111011000101001011,
    24'b001001101011000001001111,
    24'b001010101000011001000011,
    24'b000000000000000000000000,
    24'b000110110101000010010111,
    24'b000010110110000111000100,
    24'b000000110110010111010110,
    24'b000001000110011011010011,
    24'b000000010110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000100110011111010001,
    24'b000001010110011011010100,
    24'b000000010110011111001110,
    24'b000011100110001011000101,
    24'b000110010100011110001101,
    24'b000000000000000000000000,
    24'b000111110101101000101100,
    24'b001001001011000001001101,
    24'b000111111011001001010000,
    24'b001000111011000101001101,
    24'b001001111010111101001100,
    24'b001000011011000101001111,
    24'b001000011011001001001010,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001001011011000001001011,
    24'b001000001011001001010000,
    24'b001001001011000001001111,
    24'b001001111011000001010000,
    24'b000000000000000000000000,
    24'b000000010001101001000011,
    24'b000110010110010010111010,
    24'b000000110110001111000101,
    24'b000000000110011111010011,
    24'b000000000110011111001110,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000100110011111010001,
    24'b000000100110100011010010,
    24'b000001000110010011010101,
    24'b000000000110100111010000,
    24'b000010100110001111000100,
    24'b001001010110010010110100,
    24'b000000110001010000111000,
    24'b000000000000000000000000,
    24'b001010101010110101010000,
    24'b001001011010111101001100,
    24'b001000011011001001001100,
    24'b001001001011000101001011,
    24'b001000001011001001001100,
    24'b001001001011000001001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001001001011000001001111,
    24'b001000111011000101001010,
    24'b001000011011000101010000,
    24'b001000111011000101001100,
    24'b001011101001101101010000,
    24'b000000000000000000000000,
    24'b000110010100101010001010,
    24'b000001000110001011000010,
    24'b000000010110011111000100,
    24'b000000000110101011010001,
    24'b000000010110011011001110,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011111010000,
    24'b000000100110100111010000,
    24'b000001110110010111001000,
    24'b000011110110001111000010,
    24'b000100100011110001111000,
    24'b000000000000000000000000,
    24'b000101110100111100011111,
    24'b001000011010111101001010,
    24'b001000111011001001001001,
    24'b001000111011000101001101,
    24'b001000111011000101001100,
    24'b001000111011000101001111,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000011011000101001111,
    24'b001000011011001001001010,
    24'b001001001011000001001111,
    24'b001001101011000001001111,
    24'b000000000000000000000000,
    24'b000000010000111100101111,
    24'b001000000110010010110011,
    24'b000010000110101011010000,
    24'b000000100110011111000111,
    24'b000000010110100011010000,
    24'b000000110110011011010001,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010001,
    24'b000001110110011011010011,
    24'b000000000110011111010000,
    24'b000001010110011111001101,
    24'b000111000110010010110101,
    24'b000000000001011101000001,
    24'b000000000000000000000000,
    24'b001110011010010001011001,
    24'b001000101011001101001100,
    24'b001001011010111101001111,
    24'b001000011011000101001101,
    24'b001000011011001001001100,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001011,
    24'b001000111011000001010000,
    24'b001001101010111101001101,
    24'b001000000110101100101111,
    24'b000000000000000000000000,
    24'b000101100100011110001011,
    24'b000011110110000111000000,
    24'b000000110110001111010011,
    24'b000000010110011011001111,
    24'b000000010110011011010000,
    24'b000000010110010111010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110010111010110,
    24'b000000100110011111011000,
    24'b000001100110101111010001,
    24'b000100100110101011000001,
    24'b000101100100101110001110,
    24'b000000000000000000000000,
    24'b000011100011100000010011,
    24'b001001101010111101001101,
    24'b001000111010111001010001,
    24'b001000101011000101001100,
    24'b001000001011001101001011,
    24'b001000111011000001001111,
    24'b001001001011000001001111,
    24'b001000111011000101001111,
    24'b001000011011001001001101,
    24'b001000011011001001001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001010,
    24'b001000011011001001001100,
    24'b001000111011000001010000,
    24'b001001001011000001001110,
    24'b001001011011000001001010,
    24'b001001001011000101001011,
    24'b001001001011000001001100,
    24'b001001001011000001001111,
    24'b001010101010110001010001,
    24'b000000000000000000000000,
    24'b000000010001111001001111,
    24'b000110000110000110111000,
    24'b000001100110011011001110,
    24'b000001000110010111010011,
    24'b000000010110011011010001,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000010110011011010001,
    24'b000000110110010111010100,
    24'b000000010110011111010000,
    24'b000010000110010011000011,
    24'b000111010110000110111010,
    24'b000011000010011001100010,
    24'b000000000000000000000000,
    24'b000110100101100100100100,
    24'b001001101010110101001100,
    24'b001000001011000101001100,
    24'b001001011010110101010001,
    24'b001000001011001001001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001001111010111101001101,
    24'b001001001011000001001101,
    24'b001000101011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000011011001001001100,
    24'b001001001011000001001101,
    24'b001000101011001001001100,
    24'b000111111011001001001101,
    24'b001000011011001001001101,
    24'b001000011011000101001110,
    24'b000111101011001101001101,
    24'b001000111011000001001101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000110100101010010011101,
    24'b000010010110011111000111,
    24'b000001100110101111010101,
    24'b000000000110010111001111,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001101,
    24'b000000010110011111001100,
    24'b000001000110010011010010,
    24'b000000000110010011010010,
    24'b000001010110011111001111,
    24'b000100010110010111001010,
    24'b000110100101110010101001,
    24'b000000000001011100110100,
    24'b000000000000000000000000,
    24'b001111011001111101010011,
    24'b001000011011000101001101,
    24'b001000101011000101001110,
    24'b001001011011000001001101,
    24'b001001011011000001001100,
    24'b000111101011001101001100,
    24'b001001001011000001001101,
    24'b001001011011000001001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000101011000101010000,
    24'b001000101011001001001100,
    24'b001001001011001001001001,
    24'b001000111011000101001100,
    24'b001000011011000101001111,
    24'b001001001011000001001110,
    24'b001001111011001101001101,
    24'b001001110110101100111001,
    24'b000000000000000000000000,
    24'b000101010100001001111100,
    24'b000101010110010110111111,
    24'b000000100110010011001111,
    24'b000000100110011111010001,
    24'b000000100110011111010001,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010011,
    24'b000001000110010011010101,
    24'b000000010110011011010101,
    24'b000000000110010111001110,
    24'b000010000110100111001101,
    24'b000100100110001110111111,
    24'b000101110101001110010100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001101101001100101010000,
    24'b001000101011001001001011,
    24'b001000011011000101001100,
    24'b001001111010111101001100,
    24'b001000011011001101001100,
    24'b000111111011001101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001001011011000001001110,
    24'b000111111011001001001101,
    24'b001001001011000001001011,
    24'b001001101010111101001110,
    24'b001000101011001001001101,
    24'b001000011011001001001000,
    24'b001111011010000001011000,
    24'b000000000000000000000000,
    24'b000001110010101001011001,
    24'b000110000110000110110001,
    24'b000000000110011111001101,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110010111010101,
    24'b000000010110010111010100,
    24'b000000010110011111010010,
    24'b000000000110010111001101,
    24'b000001000110011011001011,
    24'b000001110110100011000010,
    24'b000100100110001011001101,
    24'b000101010100000110000011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001010011010110001001111,
    24'b000111111011000001001111,
    24'b001000101011000101001111,
    24'b001001011010110101001010,
    24'b001001001011000001001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001001011011000001001011,
    24'b001000011011001001001101,
    24'b001000011011000101001111,
    24'b001000011011000101001100,
    24'b001000101011000101010000,
    24'b001101101010001001010111,
    24'b000000000000000000000000,
    24'b000000100001110001000100,
    24'b000110010101111010101110,
    24'b000010000110011111000110,
    24'b000001000110011011001010,
    24'b000001000110010011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110100011001101,
    24'b000000000110100111001111,
    24'b000000000110011111010000,
    24'b000000110110011011010010,
    24'b000001100110010011010010,
    24'b000000000110010111010000,
    24'b000001100110011111001100,
    24'b000101000110000110111100,
    24'b000100110100000101110101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001110001010000001010000,
    24'b000111101011001001010000,
    24'b001000111011010001001111,
    24'b001000111011000101001101,
    24'b001000001011001001001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001011,
    24'b001000101011000101001110,
    24'b001001001011000001001110,
    24'b001001001011010101001011,
    24'b001101101010001001010111,
    24'b000000000000000000000000,
    24'b000000010001100101000001,
    24'b000110010101111010100100,
    24'b000010010110011011001000,
    24'b000001100110100111010100,
    24'b000000100110011111010000,
    24'b000000000110100111001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011111010101,
    24'b000000010110011111010101,
    24'b000001000110011011001110,
    24'b000001000110010011001011,
    24'b000010000110010111001100,
    24'b000101010110001010111101,
    24'b000101000011111001111001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010000001010000101011000,
    24'b000111111011010001001010,
    24'b001001011011001001001110,
    24'b001000111011001101010001,
    24'b001000111011000101001101,
    24'b001000111011000101001111,
    24'b001000001011001001001110,
    24'b001000111011000101001100,
    24'b001001001011000001001011,
    24'b001000001011001001001111,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001001001011000001001101,
    24'b001000111011000101001011,
    24'b001000011011001001001101,
    24'b001001111010111001001111,
    24'b001001001011000101001011,
    24'b001000001011001001001100,
    24'b001001101011000101001100,
    24'b001001101010111101010000,
    24'b001010100111011000111101,
    24'b000000000000000000000000,
    24'b000000000001110001000110,
    24'b000100100110000010101101,
    24'b000010110110000110111101,
    24'b000001000110010011001010,
    24'b000000000110010111001111,
    24'b000000010110100011010000,
    24'b000000000110011111001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000110110100011010100,
    24'b000000010110010111010001,
    24'b000000100110011011010010,
    24'b000011000110101011010001,
    24'b000101110110000010110101,
    24'b000101110100011110000111,
    24'b000000010001000000101011,
    24'b000000000000000000000000,
    24'b000101100101101000100001,
    24'b001010011011000101010011,
    24'b000111111011001001001111,
    24'b001000001011001001001011,
    24'b001000101011000101001011,
    24'b001000101011000101001011,
    24'b001001001011000101001011,
    24'b001000101011000101001011,
    24'b001001001011000001001011,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b000111111011001001001101,
    24'b001000011011000101001101,
    24'b001001001011000001001011,
    24'b001000011011001001001101,
    24'b001001001011000001010000,
    24'b001001011011001101001110,
    24'b001011101010110001001110,
    24'b000011100011011100010100,
    24'b000000000000000000000000,
    24'b000001100010000101010001,
    24'b000110110110000110110010,
    24'b000011010110010011000011,
    24'b000010110110011111001101,
    24'b000000010110010011010011,
    24'b000000000110011111011000,
    24'b000000000110011011010100,
    24'b000000010110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000010110100011001111,
    24'b000000000110011111001110,
    24'b000000100110011111010011,
    24'b000000110110100011010010,
    24'b000000000110011011010000,
    24'b000000100110100011010100,
    24'b000001010110010111001011,
    24'b000100010110010011000100,
    24'b000110000101000010010111,
    24'b000000010001011100111001,
    24'b000000000000000000000000,
    24'b000111110011111100100100,
    24'b001011101010101001010010,
    24'b001001001011000001001110,
    24'b001000111011000101001011,
    24'b001001101010111101001100,
    24'b001000011011000101001110,
    24'b001000111011000001001111,
    24'b001000111011000101001110,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001110,
    24'b001000111011000001010000,
    24'b001000011011001001001101,
    24'b001001001011000101001011,
    24'b001000011011000101001101,
    24'b001001001011000101001010,
    24'b001110011010010101010011,
    24'b000000000000000000000000,
    24'b000000010000110100101100,
    24'b000011000011001101110000,
    24'b000110100110011010110001,
    24'b000010010110101011001101,
    24'b000001000110011011001100,
    24'b000000010110010111010001,
    24'b000000000110011111010101,
    24'b000000010110101011011001,
    24'b000000000110010111010100,
    24'b000000000110010111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000010110011111010000,
    24'b000000010110011111001110,
    24'b000000010110011111001100,
    24'b000000100110011111001100,
    24'b000001000110010111001101,
    24'b000001010110010111001100,
    24'b000010100110010111000011,
    24'b001000100110000010101100,
    24'b000010010010101001010111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000111100101110000101101,
    24'b001010111010101001010110,
    24'b001001011011001001001100,
    24'b001000001011001001001010,
    24'b001000111010111001001100,
    24'b001000011011001101001100,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001100,
    24'b001000101011001001001101,
    24'b001000111011001001001110,
    24'b001001001011000001001100,
    24'b001100001010100101010100,
    24'b001000000101010100110000,
    24'b000000000000000000000000,
    24'b000000010001011100111011,
    24'b000101010100110110010100,
    24'b000011100110010010111110,
    24'b000001010110010011000111,
    24'b000000010110101011001000,
    24'b000000000110100011001110,
    24'b000000000110100011001111,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011001110,
    24'b000000000110011111010000,
    24'b000000010110011011001111,
    24'b000000110110011011001101,
    24'b000000110110011011001110,
    24'b000000010110011011001110,
    24'b000000010110010011001010,
    24'b000010000110011011001000,
    24'b000100100110010010111100,
    24'b000101110100111010001100,
    24'b000000000001011001000110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001011000111001000111100,
    24'b001010101010101101010010,
    24'b001010001010111101010010,
    24'b001000111010111001001110,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000001001101,
    24'b001001111010111101010000,
    24'b001100001010100001010110,
    24'b001010000101100100110001,
    24'b000000000000000000000000,
    24'b000000000000101000101011,
    24'b000001110011000001100010,
    24'b001000100101111010101100,
    24'b000011010110010111000110,
    24'b000000110110101011001000,
    24'b000000000110011111001110,
    24'b000001000110010111010011,
    24'b000000000110011111010001,
    24'b000000000110011011001111,
    24'b000000010110011011001110,
    24'b000000010110011011001101,
    24'b000000000110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011011010011,
    24'b000000010110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111010100,
    24'b000000000110011011010010,
    24'b000000000110011111010010,
    24'b000000010110100011010010,
    24'b000000000110010111001101,
    24'b000001110110010011010000,
    24'b000001000110010111001101,
    24'b000011100110010011001000,
    24'b001000010110000010110111,
    24'b000101100100001010000000,
    24'b000000010001010101000001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000010110010111000010000,
    24'b001001111000100101000011,
    24'b001100001010100001010010,
    24'b001001011010111001001101,
    24'b001000001011001001001100,
    24'b001001001011000001001101,
    24'b001000101011000101001101,
    24'b001000111011000101001100,
    24'b001000111011000101001100,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001101,
    24'b001000111011000101001100,
    24'b001001001011000101001010,
    24'b001000111011000101001011,
    24'b001000111011000101001101,
    24'b001001101010111001010010,
    24'b001101001010010101011000,
    24'b001011101000010001000111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000101100110100,
    24'b000001100010010001011110,
    24'b000110100101100010011111,
    24'b000011010101111110111000,
    24'b000010010110100011001110,
    24'b000001000110011011001101,
    24'b000001000110011111001101,
    24'b000000000110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011011010001,
    24'b000000010110011011010000,
    24'b000000010110011011001110,
    24'b000000010110011011001111,
    24'b000000000110011011010001,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000100110100111010010,
    24'b000000000110011111001111,
    24'b000000000110011111001101,
    24'b000000000110011111010000,
    24'b000000100110011011010010,
    24'b000001010110010111001100,
    24'b000010100110010011001000,
    24'b000011000110001010111110,
    24'b000111110110011110111000,
    24'b000110110100101010001010,
    24'b000001110001111001001010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001011110110001100111011,
    24'b010000111001000101011000,
    24'b001111011001010101010000,
    24'b001000101010111101001111,
    24'b001000101011000001001111,
    24'b001000101011000101001110,
    24'b001001001011000001001110,
    24'b001000101011000001001101,
    24'b001000101011000101001111,
    24'b001110011001100101011000,
    24'b010001001001001001011101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001011100111010,
    24'b000011100011011101101111,
    24'b000111000101100110100100,
    24'b000101010110010010111110,
    24'b000001100110000011000001,
    24'b000001000110001111001001,
    24'b000001010110100011001111,
    24'b000001100110100011010100,
    24'b000000110110011111010110,
    24'b000000010110011111010010,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011011001101,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000001000110010111001110,
    24'b000001000110110111010000,
    24'b000001000110110011001111,
    24'b000100010110011011001001,
    24'b000111000110001010111011,
    24'b001001110110000010101010,
    24'b000100010100011010000010,
    24'b000000000010100101010110,
    24'b000000000001000100110110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000101100101110,
    24'b000000000010001101001111,
    24'b000100100011100001110100,
    24'b000101110101001110010110,
    24'b000101110110001010111010,
    24'b000100100110011011000010,
    24'b000010110110011111001010,
    24'b000000000110001111001001,
    24'b000000000110011111001100,
    24'b000000110110011011001101,
    24'b000000110110011011001110,
    24'b000000110110011011010010,
    24'b000000110110100011010100,
    24'b000000010110011111010010,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011011010011,
    24'b000000000110011011010100,
    24'b000000000110011011010011,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000010110100111001110,
    24'b000000100110100111001101,
    24'b000001010110010011001100,
    24'b000010010110001011001101,
    24'b000011010110001011000001,
    24'b000100100110000010110110,
    24'b000110100101101110100110,
    24'b000101010101011010010111,
    24'b000101000100010110000010,
    24'b000100110011110101111000,
    24'b000100100011100101110011,
    24'b000100010011011101101100,
    24'b000100100011100101101100,
    24'b000100010011101101110000,
    24'b000101110100001101111101,
    24'b000111100100111010010101,
    24'b000110010101100110100100,
    24'b000101110101110110110000,
    24'b000100110110001010111001,
    24'b000010010110010110111111,
    24'b000010110110010011000101,
    24'b000001100110010111001101,
    24'b000000110110010111001011,
    24'b000000010110011011001100,
    24'b000000110110011011001100,
    24'b000000100110011011001101,
    24'b000000110110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011010001,
    24'b000000010110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010100,
    24'b000000000110011111010100,
    24'b000000100110010111010001,
    24'b000000010110011011010010,
    24'b000000000110011111010001,
    24'b000000000110100011010001,
    24'b000000000110011111001110,
    24'b000000100110011011001101,
    24'b000001000110011011001011,
    24'b000000100110010111001001,
    24'b000001000110010011000111,
    24'b000010010110010011000100,
    24'b000010000110100011000110,
    24'b000011010110011111000110,
    24'b000010110110011011000101,
    24'b000011000110010111000001,
    24'b000010100110010010111101,
    24'b000010110110011011000010,
    24'b000010000110010111000011,
    24'b000001000110010011000100,
    24'b000010000110010111001001,
    24'b000001110110011011001101,
    24'b000001010110011011001101,
    24'b000000100110011111001110,
    24'b000000000110100111001111,
    24'b000000010110011011001110,
    24'b000000000110011111001111,
    24'b000000000110011011010001,
    24'b000000010110011111010010,
    24'b000000100110011011010100,
    24'b000000010110011011010000,
    24'b000000010110011011001110,
    24'b000000000110011011010001,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011001111,
    24'b000000010110011011010001,
    24'b000000010110011011010001,
    24'b000000010110011111010000,
    24'b000000100110011011010001,
    24'b000000010110011011010011,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000010110100011001111,
    24'b000000100110011111001110,
    24'b000000010110011111010000,
    24'b000000100110010011001111,
    24'b000000010110011111001110,
    24'b000000010110011111001111,
    24'b000001100110010111001110,
    24'b000000110110100011001101,
    24'b000001000110100011001101,
    24'b000001000110011011001110,
    24'b000000100110011011001011,
    24'b000000110110011111001100,
    24'b000000110110011111001111,
    24'b000000100110011111010001,
    24'b000000100110100111010000,
    24'b000000010110100111001110,
    24'b000000010110011011010000,
    24'b000001000110010111010010,
    24'b000000000110011111001111,
    24'b000000000110011011010010,
    24'b000000000110011011010100,
    24'b000000010110011011010011,
    24'b000000010110011011010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011111010101,
    24'b000000100110011011010100,
    24'b000000110110010111010010,
    24'b000000110110010111010000,
    24'b000001000110011011010001,
    24'b000000010110011011010010,
    24'b000000100110011011010100,
    24'b000000010110010111010011,
    24'b000000010110011011010001,
    24'b000000000110011111001101,
    24'b000000000110100011001100,
    24'b000000000110011111001111,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010010,
    24'b000000010110011111010011,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010010,
    24'b000000010110011111010101,
    24'b000000010110011011010010,
    24'b000000010110011011001111,
    24'b000000010110011111001100,
    24'b000000000110011111001100,
    24'b000000000110011111001111,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000010110100111010010,
    24'b000000100110100111010010,
    24'b000000100110100111010010,
    24'b000000010110011111010011,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000100110100011010100,
    24'b000000000110100111010110,
    24'b000000100110011111010011,
    24'b000000010110011011010000,
    24'b000000100110100011001101,
    24'b000000010110100011001101,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000
};

assign mem_green = memory_green;

endmodule
