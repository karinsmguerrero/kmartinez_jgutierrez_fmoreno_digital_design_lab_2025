module lab2tallerdis(input logic a, b, output logic c);

endmodule 