module shift_left_nbit #(parameter N = 4) (
    input logic [N-1:0] A,
    input logic [$clog2(N):0] shift_amount,
    output logic [N-1:0] Y
);
    assign Y = A << shift_amount;
endmodule
