module lab2tallerdis_tb();

endmodule 