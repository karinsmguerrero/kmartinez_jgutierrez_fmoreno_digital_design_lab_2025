module sprite_tile(output logic [23:0] mem [0:8099]);


logic [23:0] memory [0:8099] = '{
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110100011001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011011010001,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111010001,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100011001110,
    24'b000000000110100011001110,
    24'b000000000110100011001110,
    24'b000000000110011011001101,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000000110011111001110,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000000110011111001110,
    24'b000000000110100011001110,
    24'b000000000110100011001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110100011001110,
    24'b000000000110100011001110,
    24'b000000000110011111001110,
    24'b000000010110100011001110,
    24'b000000000110011111001100,
    24'b000000000110011111001100,
    24'b000000000110011111001100,
    24'b000000000110011111001100,
    24'b000000010110011111001100,
    24'b000000010110011111001100,
    24'b000000010110011111001100,
    24'b000000000110011111001100,
    24'b000000000110011111001100,
    24'b000000000110100011001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000100110011111001110,
    24'b000000100110011111010000,
    24'b000000100110011111010001,
    24'b000000010110011011010000,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110100011010011,
    24'b000000000110100011010011,
    24'b000000000110100011010011,
    24'b000000010110100011010001,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011011010001,
    24'b000000000110011011010010,
    24'b000000000110011011010001,
    24'b000000010110100011010001,
    24'b000000010110100011010010,
    24'b000000010110100011010001,
    24'b000000010110100011010001,
    24'b000000010110100011010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000010110011011001111,
    24'b000000010110011011010000,
    24'b000000110110010111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000100110011111001101,
    24'b000000100110100011001111,
    24'b000000010110011011001111,
    24'b000000010110011011010001,
    24'b000000100110011011010011,
    24'b000000100110011011010101,
    24'b000000100110011011010101,
    24'b000000000110011111010011,
    24'b000000000110100011010010,
    24'b000000000110011111010001,
    24'b000000010110011111010001,
    24'b000000010110011111010000,
    24'b000000110110011111001111,
    24'b000001000110100011001111,
    24'b000000010110011111010000,
    24'b000000010110011111001110,
    24'b000000010110011111001100,
    24'b000000010110011111001100,
    24'b000000010110011111001100,
    24'b000000110110100111001111,
    24'b000000110110100111010010,
    24'b000001000110100111010100,
    24'b000001000110100011010011,
    24'b000000100110011011010010,
    24'b000000100110100011010100,
    24'b000000010110011111010011,
    24'b000000010110011111010011,
    24'b000000100110011111010100,
    24'b000000100110011111010100,
    24'b000000100110011111010011,
    24'b000000110110011011010011,
    24'b000001000110011011010011,
    24'b000001000110011011010011,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011011001010,
    24'b000000000110011011001011,
    24'b000000010110011011001111,
    24'b000000010110011011010001,
    24'b000000010110010111010100,
    24'b000000010110010111010101,
    24'b000000000110010011010100,
    24'b000000010110011111010010,
    24'b000000010110011011010000,
    24'b000000010110011011001111,
    24'b000000110110011111001111,
    24'b000000110110011011001100,
    24'b000001000110010111001100,
    24'b000001000110011011001011,
    24'b000001010110011111001100,
    24'b000001000110011111001011,
    24'b000000110110011011001000,
    24'b000000110110011011000101,
    24'b000001000110011011000111,
    24'b000001010110011111001011,
    24'b000001000110011011001100,
    24'b000001000110011011001101,
    24'b000001000110010111001100,
    24'b000000110110010111001101,
    24'b000000110110011011001111,
    24'b000000110110011011010000,
    24'b000000110110011011010001,
    24'b000000110110010111010011,
    24'b000000010110011011010010,
    24'b000000110110011111010001,
    24'b000001000110011011010001,
    24'b000001000110011011010001,
    24'b000001000110011011010001,
    24'b000000010110011111010001,
    24'b000000000110011011010000,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000010110100011010001,
    24'b000000000110011111001110,
    24'b000000010110011111001011,
    24'b000000000110011011001010,
    24'b000000010110011011001101,
    24'b000000110110011111010011,
    24'b000000100110011011010101,
    24'b000000100110011011010110,
    24'b000000010110010111010101,
    24'b000000100110011111010010,
    24'b000000100110011111001111,
    24'b000001000110011111001111,
    24'b000001000110011111001101,
    24'b000001100110011111001101,
    24'b000001100110011011001100,
    24'b000001010110010111001001,
    24'b000010000110010011001001,
    24'b000010000110010011001000,
    24'b000010000110010111000100,
    24'b000010000110010111000010,
    24'b000010000110010111000100,
    24'b000001110110010011000101,
    24'b000010000110010011001000,
    24'b000001100110011011001000,
    24'b000001010110011011000111,
    24'b000001010110010111001001,
    24'b000001000110011011001010,
    24'b000001000110010111001100,
    24'b000000110110011011001110,
    24'b000000110110011011001110,
    24'b000000110110011011001110,
    24'b000000110110011111001110,
    24'b000001000110011111001110,
    24'b000001000110011111001111,
    24'b000001000110011111001111,
    24'b000000010110011011001101,
    24'b000000010110011011001101,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000000110100011010000,
    24'b000000000110100011010010,
    24'b000000000110011111010001,
    24'b000000000110011111001111,
    24'b000000100110011011001110,
    24'b000000100110010111001110,
    24'b000000000110011011010100,
    24'b000000000110011011010100,
    24'b000000100110011111010101,
    24'b000000100110101111010111,
    24'b000000010110100111010010,
    24'b000001000110100111001011,
    24'b000001000110010111000010,
    24'b000010010110011011000100,
    24'b000010110110010010111101,
    24'b000101000110010110111010,
    24'b000101010101101110101011,
    24'b000110000101100010100011,
    24'b000110000101001110011101,
    24'b000101000100110010010100,
    24'b000011100100001110001000,
    24'b000010110011111010000011,
    24'b000010010011110101111111,
    24'b000010000011110101111110,
    24'b000010000011110001111110,
    24'b000100110100100010001100,
    24'b000110110101000010010110,
    24'b000110010101110010100100,
    24'b000100110101111010101000,
    24'b000100000101111110101110,
    24'b000100010110001110111000,
    24'b000011100110010110111110,
    24'b000001110110000111000010,
    24'b000010000110010011001101,
    24'b000001100110001111001011,
    24'b000001000110010111000110,
    24'b000000110110011111001111,
    24'b000000000110010111010001,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000000110100011010011,
    24'b000000000110100011010011,
    24'b000000000110100111010010,
    24'b000000100110011011001101,
    24'b000000110110011011001101,
    24'b000000000110100011010011,
    24'b000000000110101011010101,
    24'b000000000110100011010101,
    24'b000000110110010111010001,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011011010000,
    24'b000000000110100011010010,
    24'b000000000110011111010001,
    24'b000000110110011111001100,
    24'b000000110110010111001001,
    24'b000000000110010111001110,
    24'b000000000110011111010011,
    24'b000000110110011011001011,
    24'b000001110110010111001000,
    24'b000011010110011011000111,
    24'b000010100110000111000000,
    24'b000100110110011011000011,
    24'b000101100110001110111100,
    24'b000101010101110010101110,
    24'b000111000100111010001110,
    24'b000011100011101001110010,
    24'b000010000010100001010111,
    24'b000000110001101001000001,
    24'b000000000001001100110000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001001000110101,
    24'b000000010001101001000100,
    24'b000001100010101101011010,
    24'b000011010011111101110101,
    24'b000100100101000010010000,
    24'b000101100101101110100110,
    24'b000101100110000010111001,
    24'b000100010110001011000111,
    24'b000001100110001111001000,
    24'b000001010110101011010000,
    24'b000000110110100011001101,
    24'b000001000110100111001110,
    24'b000000100110011011001110,
    24'b000000010110010111010010,
    24'b000000000110011011010011,
    24'b000000000110100011001110,
    24'b000000000110100011001011,
    24'b000000000110011111001110,
    24'b000000010110011111010011,
    24'b000000010110011011010000,
    24'b000000110110011011001100,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000000110011011010010,
    24'b000000010110011011010000,
    24'b000001000110010111001011,
    24'b000001010110011011001100,
    24'b000000000110100011010010,
    24'b000000000110011111010101,
    24'b000000100110011111010000,
    24'b000011100110010111000100,
    24'b000110100101111010110001,
    24'b001000100101100010011101,
    24'b000101110100000101111100,
    24'b000010100010100001011010,
    24'b000000100001011100111111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000110001010000110000,
    24'b000010100010100001010101,
    24'b000100100100001110001000,
    24'b000110110101100110101110,
    24'b000110010110011111001000,
    24'b000011100110010111001100,
    24'b000001110110010011001011,
    24'b000001000110011011001001,
    24'b000000010110010111001001,
    24'b000000110110011011001110,
    24'b000000100110011111001001,
    24'b000000100110011111001000,
    24'b000000100110011011001011,
    24'b000000010110010011001111,
    24'b000000100110011011010001,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011001111,
    24'b000000100110011011001101,
    24'b000000000110011011010010,
    24'b000000000110100011011010,
    24'b000000000110011111010111,
    24'b000001010110010111001111,
    24'b000011010110010011001001,
    24'b000101110110001111000000,
    24'b000101110101000110011111,
    24'b000001100010101101100011,
    24'b000000100001000000110101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010000100011100100110101,
    24'b011010100110001001011110,
    24'b100001000111101001111001,
    24'b100100101000011110000110,
    24'b101000111001100110010111,
    24'b101010011001111010011100,
    24'b101001101001101110011001,
    24'b101000011001011010010101,
    24'b100100111000100010001000,
    24'b100000100111011101110111,
    24'b011000000101101101010111,
    24'b001110000011100100110100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000100001011101000001,
    24'b000010000011000001110001,
    24'b000111000101010010100100,
    24'b000110000110010010111110,
    24'b000010000110010011000011,
    24'b000000100110100111001010,
    24'b000000100110100111001000,
    24'b000001100110001111001000,
    24'b000001010110001111001011,
    24'b000000110110101011010010,
    24'b000000000110101111010110,
    24'b000000000110100111010101,
    24'b000000000110010111010100,
    24'b000000010110011011010001,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110101011001110,
    24'b000000110110011011001000,
    24'b000000010110011011010000,
    24'b000000000110100111011100,
    24'b000000100110010011010011,
    24'b000110100110010111000000,
    24'b000111000100110110010010,
    24'b000001110010010101010001,
    24'b000000000000100100101001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010111000101000001010000,
    24'b101001001001011010010101,
    24'b110101111100100111000011,
    24'b111011111110000011010111,
    24'b111100111110001111010111,
    24'b111100011110000111010010,
    24'b111100111110001111010011,
    24'b111100001110000011010011,
    24'b111100101110000111011001,
    24'b111100101110000111011001,
    24'b111100101110000111011001,
    24'b111100011110000011011001,
    24'b111100101110000111011010,
    24'b111100111110001011011011,
    24'b111011111110010011010111,
    24'b111011111110010111011010,
    24'b111010111110000111011011,
    24'b110010011100001010111111,
    24'b100101101001000110001110,
    24'b010010100100100001001000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000001100010111001100010,
    24'b000101100101010010100001,
    24'b000011100110000010111100,
    24'b000000110110011111000101,
    24'b000000110110011011001101,
    24'b000000000110011011010011,
    24'b000000010110011011010100,
    24'b000000110110100111010100,
    24'b000000100110011011010000,
    24'b000001000110010111001110,
    24'b000000110110010111010000,
    24'b000001000110011011010001,
    24'b000000100110011111010001,
    24'b000000010110011011010000,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000010110011111001101,
    24'b000001110110011011001001,
    24'b000011100110011011000110,
    24'b000100010110001010111101,
    24'b000101000101011010100000,
    24'b000001100010110101100011,
    24'b000000000001001000110010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010110100101000101001111,
    24'b101011101010010010100100,
    24'b111001111101101111011010,
    24'b111011111110001011011010,
    24'b111011101110001011011010,
    24'b111011001101111011010110,
    24'b111101001110011011011110,
    24'b111100101110010011011100,
    24'b111101011110010111011110,
    24'b111011011101110111011000,
    24'b111100011110001111010100,
    24'b111011111110000111010010,
    24'b111100011110001011010101,
    24'b111100001110000111010101,
    24'b111100001110001011010110,
    24'b111100011110001011010110,
    24'b111100011110001011010110,
    24'b111100001110000011010110,
    24'b111101111110010111100000,
    24'b111100011110001011011111,
    24'b111011101110000111011101,
    24'b111011111110011011011101,
    24'b111011011110011111011010,
    24'b110110111101011011001001,
    24'b101011011010100110011110,
    24'b010011000100100001000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000111100110010,
    24'b000010110011000101100011,
    24'b000100010101101010100111,
    24'b000011000110100011000000,
    24'b000001000110101011001111,
    24'b000001100110011011010010,
    24'b000010100110000111001011,
    24'b000010010110001011000110,
    24'b000001000110011011000110,
    24'b000000110110010111001101,
    24'b000000110110011011001110,
    24'b000000110110011011001110,
    24'b000000010110011011010000,
    24'b000000010110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000001010110010111010001,
    24'b000010100110011011001101,
    24'b000101100101110110110011,
    24'b000100000011100101110000,
    24'b000000100001000100101011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001010000010000100100001,
    24'b100010100111111101111010,
    24'b110101011100101111000010,
    24'b111010001101111011010111,
    24'b111010111110000011010111,
    24'b111100001110001011011010,
    24'b111011101110000111010111,
    24'b111100011110010011011010,
    24'b111011011101111111010110,
    24'b111100111110010011011011,
    24'b111101001110010011011011,
    24'b111011111101111011010101,
    24'b111100111110001011011000,
    24'b111100001101111111010000,
    24'b111100011110000111010010,
    24'b111100111110000111010101,
    24'b111100111110000111010110,
    24'b111100111110000111010110,
    24'b111100111110001011010111,
    24'b111100111110000111010101,
    24'b111100011110001011010110,
    24'b111011111110000011011000,
    24'b111011111110000011011011,
    24'b111100111110010011011111,
    24'b111100001110000111011000,
    24'b111100001110001111010101,
    24'b111011101110001011010011,
    24'b111100101110010011011000,
    24'b111100011110001011011010,
    24'b110100001100011111000010,
    24'b011110010111010001110001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001100000111011,
    24'b000011100100000001111101,
    24'b000101110110000010110110,
    24'b000011100110010111001011,
    24'b000001110110010111010000,
    24'b000000110110011011010000,
    24'b000000010110100011010010,
    24'b000001000110010111001110,
    24'b000001000110010111001110,
    24'b000000110110011011001110,
    24'b000000110110011011010000,
    24'b000000100110011111010001,
    24'b000000000110011111010001,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000010110011011001111,
    24'b000000010110011011001111,
    24'b000000000110010111001110,
    24'b000000000110011011010000,
    24'b000000000110011111010001,
    24'b000000000110011111010100,
    24'b000000000110011111010000,
    24'b000000010110011011001111,
    24'b000000000110011111010100,
    24'b000000000110011111010011,
    24'b000000100110010011001100,
    24'b000001010110101011010100,
    24'b000001000110100011001111,
    24'b000100000110010010111101,
    24'b000110100101010110100101,
    24'b000001000010000101010110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100100001000001001111101,
    24'b111000001101000011001011,
    24'b111101001110001111011100,
    24'b111011111110001011011001,
    24'b111011111110001011011001,
    24'b111011111110001111011001,
    24'b111100001110001011010111,
    24'b111100101110000111011000,
    24'b111100101110000111011000,
    24'b111100111110001011011000,
    24'b111100101110000011010110,
    24'b111100111110001011010101,
    24'b111100111110000111010100,
    24'b111101001110000111010100,
    24'b111100011110000011010110,
    24'b111100101110000111011000,
    24'b111100101110000111011000,
    24'b111100101110000111011001,
    24'b111100101110000111011001,
    24'b111100101110000111011001,
    24'b111100101110000011010111,
    24'b111100101110000111010111,
    24'b111100011110000111010110,
    24'b111100011110000111011000,
    24'b111100011110000011011001,
    24'b111100101110000111011000,
    24'b111100011110001111011000,
    24'b111100011110001111011010,
    24'b111100101110000011011010,
    24'b111101011110000011011111,
    24'b111100101110000111011011,
    24'b111011011110000111010110,
    24'b110111111101010111001000,
    24'b011111110111010101101110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000010000010010101010111,
    24'b000111010101101110101001,
    24'b000011100110100011001011,
    24'b000000010110010111010001,
    24'b000001000110101011010101,
    24'b000000110110100111010010,
    24'b000000000110011011010000,
    24'b000000000110011011010000,
    24'b000000010110011011010010,
    24'b000001000110011111010001,
    24'b000000010110011011001111,
    24'b000000010110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000010110011011010000,
    24'b000000000110011011010011,
    24'b000000000110011111010011,
    24'b000000010110011011001110,
    24'b000000010110011111001100,
    24'b000000000110011111010001,
    24'b000000000110011011010011,
    24'b000000000110010111001111,
    24'b000010100110100011001010,
    24'b000100100110001110111100,
    24'b000100100100110010001101,
    24'b000000000001000000110001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010111000101100001011010,
    24'b110111111101001111001011,
    24'b111100111110001011011000,
    24'b111100011101111111010110,
    24'b111100001101111111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000111011010,
    24'b111100111110001011100001,
    24'b111100111110000011011011,
    24'b111100101110000011010100,
    24'b111110001110100011011011,
    24'b111100011110001111011001,
    24'b110111101101010011001111,
    24'b010101010100111101001100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001110101001001,
    24'b000101000100111010010011,
    24'b000101110110011110111110,
    24'b000010010110011011001001,
    24'b000000010110110011010111,
    24'b000000100110100111010011,
    24'b000000110110011011001110,
    24'b000001000110010111001100,
    24'b000001000110100011010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000100110011111001111,
    24'b000000010110011011010000,
    24'b000000000110011011010001,
    24'b000000100110011011001101,
    24'b000000000110011111001110,
    24'b000000010110011011001110,
    24'b000000100110011011001011,
    24'b000000000110011011001110,
    24'b000000110110100011001101,
    24'b000110110110011110110110,
    24'b000011100011101101110000,
    24'b000000000001000000110000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101100111010110110110001,
    24'b111010101110000011011101,
    24'b111101001110001111011010,
    24'b111101111110011011011100,
    24'b111100101110000111010111,
    24'b111100111110001011011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000111010111,
    24'b111100001110000111011001,
    24'b111100111110001111011010,
    24'b111100101110000011010110,
    24'b111100101110000111010110,
    24'b111011101110000011010111,
    24'b111010111110000011010110,
    24'b111011101110010011011011,
    24'b101000111001010110001101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010000111100101010,
    24'b000100010011111001110101,
    24'b000101110110010010110110,
    24'b000000010110100011001111,
    24'b000001110110100011010001,
    24'b000010010110000011001001,
    24'b000010000110011011001101,
    24'b000000010110100111001111,
    24'b000000000110011111001111,
    24'b000001000110011111001111,
    24'b000000010110011011001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000010110011011001111,
    24'b000000010110011011010000,
    24'b000000100110011111010001,
    24'b000000110110011011001110,
    24'b000000000110011011010010,
    24'b000000000110011111010010,
    24'b000000100110011011001101,
    24'b000001110110000111000001,
    24'b000110110110010010110100,
    24'b000001110011000001100101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010101010100010101000110,
    24'b110111111101010011001010,
    24'b111010101110001011010010,
    24'b111100101110001111011010,
    24'b111100001101101111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000011010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000111010111,
    24'b111011111110001011010101,
    24'b111100111110001111011001,
    24'b111100001101110111010110,
    24'b111100101101111111011000,
    24'b111101011110010011011100,
    24'b111011011101111111010011,
    24'b111011101110000011010010,
    24'b111101111110010111010111,
    24'b110010111100011111000001,
    24'b010000110100001000111110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000110100101000,
    24'b000011000011100101110000,
    24'b000100110110010010110110,
    24'b000010110110000011000011,
    24'b000010010110010011010011,
    24'b000000000110010011010001,
    24'b000000000110101111010000,
    24'b000000000110100011001101,
    24'b000001000110011011010001,
    24'b000000010110011011001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011001111,
    24'b000000010110011011010000,
    24'b000000110110100011010000,
    24'b000000100110011111010011,
    24'b000000010110011011010100,
    24'b000001000110100111010111,
    24'b000010000110011111001110,
    24'b000111110110000010101111,
    24'b000010110010101001011000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b011111010111010001101111,
    24'b111001101101100111010011,
    24'b111011011110001111011100,
    24'b111011101110001111011011,
    24'b111100111110001011011001,
    24'b111100111110000011010100,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000111010110,
    24'b111100001110001011010100,
    24'b111100011110000111010110,
    24'b111100101110000111011001,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100101110001011010011,
    24'b111100101110010011010100,
    24'b111010111110001111011010,
    24'b111000001101111011010111,
    24'b011000000101110001010111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000100010011101001101100,
    24'b000111010110000110110010,
    24'b000000110110001011001111,
    24'b000000000110100111011011,
    24'b000000010110101011010011,
    24'b000000100110011011001011,
    24'b000000100110011011010010,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010010,
    24'b000000000110011111010000,
    24'b000000110110100011010001,
    24'b000000110110011011001110,
    24'b000000000110010111010001,
    24'b000001010110100011010001,
    24'b000010100110001111001001,
    24'b000101110110000010110110,
    24'b000010110011000101100101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100100111000111110001011,
    24'b111000101101101011010001,
    24'b111101101110101011100000,
    24'b111010101101110111010110,
    24'b111100001110001011011100,
    24'b111100011110000111010111,
    24'b111101011110001011010100,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010110,
    24'b111100101110001011010101,
    24'b111100101110000111010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100011110001011010110,
    24'b111011011110000111010101,
    24'b111100111110011111011110,
    24'b111010011110000111011001,
    24'b111010001110010011100010,
    24'b100000000111111010000001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000011010011100001101101,
    24'b000100100110011110111101,
    24'b000000100110011111001111,
    24'b000001100110011111010001,
    24'b000001010110010111001110,
    24'b000000010110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010010,
    24'b000000000110011111010010,
    24'b000000010110011111010011,
    24'b000001000110100111010010,
    24'b000001010110011111001110,
    24'b000000100110011111001101,
    24'b000001110110011011000101,
    24'b000110010110001110110011,
    24'b000011110011100001101111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100110111001010110001110,
    24'b111010111110000011010100,
    24'b111101011110010011011111,
    24'b111100101101111111011001,
    24'b111101011110001111010110,
    24'b111101001110010011010100,
    24'b111011111110000111010101,
    24'b111100001110000111011010,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100011110001111011011,
    24'b111011101101110111010101,
    24'b111011111101110011010101,
    24'b111011111101111111011010,
    24'b111011111110001111100001,
    24'b100100011000011110000110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000011010100010101110110,
    24'b000111010110100110111101,
    24'b000011000110001011001101,
    24'b000001100110010011010101,
    24'b000000100110100111010010,
    24'b000000100110100011010100,
    24'b000000010110011011010011,
    24'b000000000110011011010010,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010010,
    24'b000000000110011111001111,
    24'b000000000110011011010001,
    24'b000000000110011111010101,
    24'b000000000110011011010010,
    24'b000001100110011111001101,
    24'b000001000110011111001111,
    24'b000000110110011011001011,
    24'b000100000110001110111100,
    24'b000101000100100010000001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100101101001010010001101,
    24'b111010111110000111010001,
    24'b111100101110001011010011,
    24'b111011111101110011010000,
    24'b111100111101111011010011,
    24'b111101011110001011010011,
    24'b111100101110001011010011,
    24'b111100011110001011011000,
    24'b111100011110001011011010,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000011011000,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110000111010110,
    24'b111100101110000111011000,
    24'b111100101110000111011000,
    24'b111011111110000111010101,
    24'b111100111110001011011001,
    24'b111101111110001011011010,
    24'b111101001101110111010100,
    24'b111100011101110011010110,
    24'b111011011101111011011000,
    24'b100001010111101101111001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000111010100111110001011,
    24'b000100100101111111000011,
    24'b000001000110010111010000,
    24'b000000100110011111010000,
    24'b000000110110100011010100,
    24'b000000000110011111010101,
    24'b000000000110011111010110,
    24'b000000000110100011010100,
    24'b000000000110011111001101,
    24'b000000000110011111001011,
    24'b000000000110011111001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100011010011,
    24'b000000010110011011001101,
    24'b000000100110011011001110,
    24'b000000000110011111010101,
    24'b000000010110011111010011,
    24'b000010100110100111001110,
    24'b000000110110010111001011,
    24'b000010100110010111000111,
    24'b000101100101010010011111,
    24'b000000000000111100110011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100001110111111101111001,
    24'b111010011110000011010110,
    24'b111011101110000111010010,
    24'b111100001110000011010001,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100101110001011010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111101001110000111011010,
    24'b111100101101111111011000,
    24'b111100001101110111010111,
    24'b011001110101110101100000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000110001100001000000,
    24'b000110110101100110100110,
    24'b000010100110100111000100,
    24'b000001100110011111001110,
    24'b000001000110010011001110,
    24'b000000110110100011010111,
    24'b000000000110011011011000,
    24'b000000010110100011010101,
    24'b000000010110100011001011,
    24'b000000000110011111001010,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001101,
    24'b000000000110011111001011,
    24'b000000000110011111001110,
    24'b000000110110100011010100,
    24'b000000100110010011001010,
    24'b000001100110001110111101,
    24'b000110100110000010100101,
    24'b000000010010000001001100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b011001110101101001010101,
    24'b111010001101101111011000,
    24'b111100001110000111011010,
    24'b111011111101110111010011,
    24'b111100101110001011010100,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010110,
    24'b111100001110001011010111,
    24'b111100011110000111010111,
    24'b111100001101111111010101,
    24'b111101011110001111011010,
    24'b111101001110001011011010,
    24'b111100111110001011011010,
    24'b111011101101111111010110,
    24'b001111110011100100110011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000110010011001010010,
    24'b000101110110000010110011,
    24'b000011000110010111000011,
    24'b000001100110001011001011,
    24'b000001010110010111010010,
    24'b000000100110011011010001,
    24'b000000100110010111010000,
    24'b000000100110010111010001,
    24'b000000010110011011010001,
    24'b000000000110011111010101,
    24'b000000000110011111010011,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000110110010111010000,
    24'b000000000110100011010000,
    24'b000000000110100111001011,
    24'b000000110110011011001100,
    24'b000000010110001111010010,
    24'b000001010110010011001111,
    24'b000101100110010110110100,
    24'b000001110011001001011100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001101100010011100100000,
    24'b111001111101100011010001,
    24'b111101001110011111100010,
    24'b111100101110000111011001,
    24'b111100101110000011010100,
    24'b111100011110000111010100,
    24'b111100011110000011010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111101001110010111011010,
    24'b111011011101111111010100,
    24'b111100001110000111010111,
    24'b111101001110010111011010,
    24'b111100001101111011001101,
    24'b111001001101100011010011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000011010011111001111011,
    24'b000011010101110110110010,
    24'b000001010110000111001111,
    24'b000001010110011011010010,
    24'b000001000110100111001111,
    24'b000000110110011011001110,
    24'b000001000110010011010010,
    24'b000000100110010011010101,
    24'b000000000110011011010100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000001010110011111010100,
    24'b000000000110011111010100,
    24'b000000000110011011010000,
    24'b000001000110011011001111,
    24'b000001100110010011010100,
    24'b000011010110000111000110,
    24'b000101010101000110010010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110010101011111010110101,
    24'b111100001110010111011100,
    24'b111011001110000011011000,
    24'b111100111110001111011000,
    24'b111100101110000011010100,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010110,
    24'b111100111110001011010010,
    24'b111100101110010011100000,
    24'b101101011010100110101100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001000100101101,
    24'b000110110101101010100100,
    24'b000001000110000111001010,
    24'b000000010110011011010010,
    24'b000000010110100011010000,
    24'b000000010110011011010000,
    24'b000001000110011011010001,
    24'b000000100110010111010001,
    24'b000000000110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000000110011011010011,
    24'b000000010110010111010100,
    24'b000000110110010011010011,
    24'b000010010110001111001100,
    24'b000111100110001010110100,
    24'b000001010010010101010111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100000110111100101110111,
    24'b111011111110010011011110,
    24'b111010111110001011011001,
    24'b111011011110001011011001,
    24'b111100001110000111010100,
    24'b111100111110001011010110,
    24'b111100101110000111011001,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010110,
    24'b111011111110000011010011,
    24'b111100101110000111011101,
    24'b111011111110010011011110,
    24'b011001000101100101011001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000001110010111001100000,
    24'b000011110110010010111011,
    24'b000001010110011111001100,
    24'b000000000110011011010010,
    24'b000000000110011111010011,
    24'b000000100110011111001110,
    24'b000000110110011011001011,
    24'b000000010110011011001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100111001101,
    24'b000000110110010111001101,
    24'b000001010110010011010100,
    24'b000000110110010011010101,
    24'b000011010110010110111111,
    24'b000101010100100010000000,
    24'b000000000000111000101110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111000111101100111010111,
    24'b111011001110000111011011,
    24'b111011011110000011011000,
    24'b111100011110001011011001,
    24'b111100101110000011010110,
    24'b111100111110000011011000,
    24'b111100101110000111011001,
    24'b111100101110000111011001,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000011011001,
    24'b111100111110000011011001,
    24'b111100111110000011011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100011110001011010101,
    24'b111100011110001111010111,
    24'b111101001110000111011000,
    24'b111011101101111011010101,
    24'b110110111101011011001111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000100110101011110010010,
    24'b000100000110010110111110,
    24'b000001000110010011010010,
    24'b000000000110011011010100,
    24'b000000000110101011001100,
    24'b000000000110100011001000,
    24'b000000010110011011010001,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011011010010,
    24'b000000000110101111001011,
    24'b000000110110010111001000,
    24'b000001110110001011010001,
    24'b000001010110011011010101,
    24'b000100000110000010101101,
    24'b000000000001100000111011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101100101010110110101001,
    24'b111011011110010011011101,
    24'b111011101110000111011001,
    24'b111100011110001111011010,
    24'b111100111110000111011000,
    24'b111101001110000011011001,
    24'b111100111110000011011001,
    24'b111100101110000111011001,
    24'b111100101110000111011001,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000011011001,
    24'b111100111110000011011001,
    24'b111100111110000011011000,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100011110001011010111,
    24'b111101101110001011010110,
    24'b111011111101111011010110,
    24'b111010011110010011011001,
    24'b100011001000001110000100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000110010011001001010,
    24'b000111100110011010110100,
    24'b000010000110000111001111,
    24'b000000100110001111010011,
    24'b000000100110101011001101,
    24'b000000000110100111001101,
    24'b000000000110010111010101,
    24'b000000000110011011010100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001100,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110100011001110,
    24'b000000000110100011001100,
    24'b000000100110011111010000,
    24'b000000110110010011011000,
    24'b000000000110100011001111,
    24'b000001000110100111001011,
    24'b000001100110011011001111,
    24'b000011010110001011000110,
    24'b000101010100101010001000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001100000010110000101001,
    24'b111101001110100111100101,
    24'b111100111110010011011100,
    24'b111100001101111111010110,
    24'b111100001110001011010111,
    24'b111100001110001011010101,
    24'b111100101110001011010101,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000111010100,
    24'b111100101110010011011011,
    24'b111011101110000111011011,
    24'b111011101110000011011001,
    24'b111001101101100011010010,
    24'b001010000001111100011011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000100100101000110001111,
    24'b000010110110011011001001,
    24'b000010110110001011001100,
    24'b000001110110101011010010,
    24'b000000000110100011010111,
    24'b000000000110100011001111,
    24'b000000000110011111001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001100,
    24'b000000000110011111001111,
    24'b000000000110011011010010,
    24'b000000000110011111001111,
    24'b000000000110011111001100,
    24'b000000010110011111010000,
    24'b000000110110010011010110,
    24'b000000100110011011001101,
    24'b000000100110101111000111,
    24'b000010100110101011001101,
    24'b000111010110001010111010,
    24'b000001000010010101010000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101101111010111110101010,
    24'b111011001101111111010111,
    24'b111100011110000011011000,
    24'b111100111110001011011000,
    24'b111100001110001011010101,
    24'b111011111110001111010101,
    24'b111100001110001011010101,
    24'b111100101110000111010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110001111010110,
    24'b111011101110000011010111,
    24'b111100011110010011011100,
    24'b111100011110001011011011,
    24'b111011111110000111011010,
    24'b100100011000100010000010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000001010010011001010111,
    24'b000110110110011010111101,
    24'b000010010110000011001000,
    24'b000001010110010111001111,
    24'b000000000110011011010010,
    24'b000000000110011111001101,
    24'b000000000110011111001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000010110011011010001,
    24'b000000110110010111010100,
    24'b000001100110010011001101,
    24'b000000000110110011000101,
    24'b000010000110011111000100,
    24'b000111010100110110011001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001011000010100000101000,
    24'b111001011101101111010100,
    24'b111101101110100011011110,
    24'b111101101110001111011000,
    24'b111100101110000111010100,
    24'b111100011110001011010101,
    24'b111011111110001111010101,
    24'b111100001110001011010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111011111110000111011000,
    24'b111011101110000011011000,
    24'b111100001110000011011001,
    24'b111100001110000011011000,
    24'b111010011101111111011001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000111000101111,
    24'b000111110101100010011111,
    24'b000010110110010111001010,
    24'b000001110110001111010001,
    24'b000001000110011011001110,
    24'b000000000110011011001100,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000010110011011010010,
    24'b000000110110010111010010,
    24'b000001010110010011001111,
    24'b000000000110110011001000,
    24'b000011110110100111000000,
    24'b000001110010100001100100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100010101000011110001000,
    24'b111010111110000111011001,
    24'b111011111101111111010010,
    24'b111101001110000011010101,
    24'b111100111110000011010011,
    24'b111100011110001011010101,
    24'b111011111110001111010101,
    24'b111100001110001011010111,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100011110001111011000,
    24'b111100001110000111011001,
    24'b111100101110000111011001,
    24'b111101001110001111011011,
    24'b111011101110000111011010,
    24'b011010100110001101011111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000110000100000101111000,
    24'b000010010110001011000000,
    24'b000001100110010011010101,
    24'b000000110110011011001110,
    24'b000000000110011111001111,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011011010100,
    24'b000000010110011011010010,
    24'b000000110110011011001110,
    24'b000001000110011011001111,
    24'b000000010110101011001011,
    24'b000100110110001010101101,
    24'b000000100001001000111011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110111011101100011010111,
    24'b111100001110010011011110,
    24'b111100111110001111011000,
    24'b111101001110000011010101,
    24'b111101001110000011010101,
    24'b111100101110001011010101,
    24'b111100001110001011010111,
    24'b111100101110000111010111,
    24'b111100101110000011011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100101110000111010111,
    24'b111100001110001011011001,
    24'b111100111110001011011001,
    24'b111100011101111111010100,
    24'b111011101101111111010111,
    24'b110111101101010111010000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001111101001011,
    24'b000101100110011010111010,
    24'b000001100110010111010001,
    24'b000000010110011011010000,
    24'b000000000110011111010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010011,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010010,
    24'b000000000110011011010101,
    24'b000000010110011011010010,
    24'b000000110110011011001100,
    24'b000000100110100011001100,
    24'b000010110110011111001101,
    24'b000101010101001010010010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001101100011011000101111,
    24'b111100001110011011011110,
    24'b111100111110010011011110,
    24'b111100111110010111011100,
    24'b111100111110000111010111,
    24'b111101001110000011010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000011011001,
    24'b111100111110000011011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000011010101,
    24'b111101011110001011010110,
    24'b111100101110001111011010,
    24'b111100111110101011100101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000110100101110,
    24'b000111110101110010100101,
    24'b000010100110100011001010,
    24'b000000100110011111010001,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111001110,
    24'b000000000110011111001101,
    24'b000000000110011111010010,
    24'b000000000110011011010110,
    24'b000000010110011011010011,
    24'b000000110110011011001011,
    24'b000000010110100011001000,
    24'b000011110110001011001000,
    24'b000011010011101001101111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100101011001000110001010,
    24'b111101011110001111010110,
    24'b111100001110000011011010,
    24'b111011011110000111011001,
    24'b111100111110000011011001,
    24'b111100111101111111010110,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000011011001,
    24'b111100111110000011011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111101001110000111010111,
    24'b111100111110000011010101,
    24'b111100001110000111011000,
    24'b111011101110001011011100,
    24'b100001010111100101110100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000110010100011010000011,
    24'b000010110110010110111110,
    24'b000000110110010111001110,
    24'b000000100110011011001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010010,
    24'b000000010110011011010011,
    24'b000000010110011011010000,
    24'b000000010110011011001110,
    24'b000000010110011111001111,
    24'b000100110110010110111011,
    24'b000001100010001101000110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110110011101001011001101,
    24'b111101011110010011011001,
    24'b111011111110001011011000,
    24'b111011111110001111011000,
    24'b111100011110000011010110,
    24'b111101001110001011011000,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000011010111,
    24'b111100101110001011011001,
    24'b111010111101101011010010,
    24'b111100001110000011011000,
    24'b110001101011111010111010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000001110010110001011011,
    24'b000011110101111110110010,
    24'b000001000110011111001101,
    24'b000000100110011111010110,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011011010000,
    24'b000000010110011011001110,
    24'b000000100110011111001110,
    24'b000101010110001010110001,
    24'b000000000001000100110001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111010011110000011011001,
    24'b111011101101110011010000,
    24'b111101011110011011011100,
    24'b111011011110000111010101,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000011011000,
    24'b111011101101110111010110,
    24'b111100101110000111011001,
    24'b111010011101111111011010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001100001000001,
    24'b000110010110011010110011,
    24'b000001000110011111001011,
    24'b000000000110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110011011010001,
    24'b000000010110011011010000,
    24'b000000010110011011001110,
    24'b000001100110100011001100,
    24'b000100100101010110011100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001100010010110000101001,
    24'b111010111101111111010101,
    24'b111101001110001011010101,
    24'b111100001110000111010101,
    24'b111011101110000011010101,
    24'b111100111110001011011000,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111011001,
    24'b111101101110010011011100,
    24'b111100011110001011011011,
    24'b001101100010101000100101,
    24'b000000000000000000000000,
    24'b000000000000111000110001,
    24'b000111110110010010101100,
    24'b000001000110011011001001,
    24'b000000000110011011010000,
    24'b000000010110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000100110011111010001,
    24'b000001010110001011000100,
    24'b000101100100101010001000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100000100111100101110110,
    24'b111100101110001111011001,
    24'b111101011110001011010110,
    24'b111100001101111011010100,
    24'b111100101110010011011001,
    24'b111100011110000011010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110001011011010,
    24'b111100001101111111010111,
    24'b111100111110001011011010,
    24'b111101101110001111011011,
    24'b011010110101110001010111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001000100101110110011111,
    24'b000001110110010111000111,
    24'b000000000110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111001111,
    24'b000000010110011011001111,
    24'b000000010110011011010000,
    24'b000001000110100111010100,
    24'b000011000110010011000100,
    24'b000101100011110001110011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101111011011001010101100,
    24'b111101001110001011010111,
    24'b111101001110001011011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110001011010111,
    24'b111100011110001011010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111011001,
    24'b111100011110000011011000,
    24'b111101101110000111011000,
    24'b100101011000100110000011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000111010100111110001100,
    24'b000010010110010011000110,
    24'b000000000110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011011001111,
    24'b000000010110011011010001,
    24'b000001000110100111010101,
    24'b000011110110010111000100,
    24'b000100100011000001011111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111010111110000011011001,
    24'b111100101110000011010100,
    24'b111100111110001011011010,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100011110000011011000,
    24'b111100011110000011011000,
    24'b111110001110001011010111,
    24'b101011001010001110011110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000100000011101101110101,
    24'b000010100110010011000110,
    24'b000000000110011111001101,
    24'b000000000110011111001110,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011011001111,
    24'b000000010110011011010001,
    24'b000001000110100111010101,
    24'b000011110110010011000011,
    24'b000011010010100001010100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111010011101111011010101,
    24'b111101001110001011010111,
    24'b111100011110000111011010,
    24'b111100111110000011011001,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100011110000011011000,
    24'b111100011110000011011000,
    24'b111110011110010011011001,
    24'b101110011011001110101101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000001010010101101100010,
    24'b000011000110010011000110,
    24'b000000000110011111001111,
    24'b000000010110011011001111,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111001111,
    24'b000000110110011011001110,
    24'b000000010110001111001110,
    24'b000100000110010011000011,
    24'b000001010010001001001101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111001011101101111010010,
    24'b111101001110010011011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100011110001011010111,
    24'b111100001110001011010111,
    24'b111100101110000011011000,
    24'b110010011100001110111010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000100010011001011000,
    24'b000011010110010110111111,
    24'b000000100110010111010000,
    24'b000000100110010111010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010000,
    24'b000000110110010111010000,
    24'b000000010110001111001110,
    24'b000011100110001011000000,
    24'b000001000010000001001011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111010001101111111010110,
    24'b111100101110001011010110,
    24'b111100101110001011010111,
    24'b111100101110000111010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100001110000111010111,
    24'b111011111110001111010111,
    24'b111100111110001011011010,
    24'b110100111100110111000011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000100010010001010100,
    24'b000011000110010110111100,
    24'b000000100110010111010001,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010000,
    24'b000000110110010111010001,
    24'b000000010110001111010000,
    24'b000011110110000111000000,
    24'b000001000001111001001001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111010101101111111011001,
    24'b111100111110000111010111,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100001110000111010111,
    24'b111011111110001111010111,
    24'b111011111110001011011001,
    24'b110100101100110111000011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000100010000101010110,
    24'b000011100110010010111011,
    24'b000000000110011011001111,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000010110011111010001,
    24'b000000110110010111010010,
    24'b000000010110001111010000,
    24'b000011110110001111000001,
    24'b000000110001111101001010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111010011101111011010111,
    24'b111101001110001011011001,
    24'b111100101110000111011001,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100011110001011010111,
    24'b111011111110001111010111,
    24'b111100001110001011010111,
    24'b110010111100011010111011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000100010001001011001,
    24'b000011000110010010111101,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000100110100011010010,
    24'b000000110110010111010010,
    24'b000001010110011111010100,
    24'b000100010110011011000100,
    24'b000001110010010101010000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111011101110000111011011,
    24'b111101001110000111011000,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100011110000011010110,
    24'b111100011110001111011000,
    24'b111011101110001011010110,
    24'b111100001110001011010111,
    24'b110001001011111110110101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000001100010101101100100,
    24'b000011000110010010111111,
    24'b000000000110100011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010001,
    24'b000001000110011011010010,
    24'b000001000110011011010010,
    24'b000011000110011011000100,
    24'b000011000010111001011011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111001111101101111010101,
    24'b111100101110000011010110,
    24'b111100011110000011010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111011111110001111010111,
    24'b111100101110000111011000,
    24'b101101011010111110101000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000011010011011101110011,
    24'b000010100110010111000010,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000010110011111010000,
    24'b000001010110100011010010,
    24'b000000110110010111001111,
    24'b000010000110011111000110,
    24'b000101000011101101101001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110101101100101011000100,
    24'b111101001110000111010110,
    24'b111100101110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110001011011000,
    24'b111100001110000111010110,
    24'b111100001110001111011000,
    24'b111101001110000011011001,
    24'b100111101001101010010100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000101100100010010000010,
    24'b000010010110011111000100,
    24'b000000000110011111010011,
    24'b000000000110011111010001,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111010001,
    24'b000000010110011111001111,
    24'b000000100110100011001110,
    24'b000000100110010111001100,
    24'b000000110110011011000111,
    24'b000101000100010001111011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101010111010000110011011,
    24'b111101001110010111011001,
    24'b111100101110000111010011,
    24'b111100001110000111010110,
    24'b111100001110001011011000,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000011010110,
    24'b111100101110000111011000,
    24'b111011111101111011010110,
    24'b111100011110000111011000,
    24'b111011111110000111010111,
    24'b100000000111101001111000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001000000101010110011111,
    24'b000001010110010111001000,
    24'b000000000110011111001100,
    24'b000000000110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111010001,
    24'b000000000110011111001111,
    24'b000000010110011111001101,
    24'b000000100110010111001010,
    24'b000000100110010111001100,
    24'b000101110100111110010001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010101010100110101001010,
    24'b111011111110000111010111,
    24'b111100011110001011010101,
    24'b111100001110001011011000,
    24'b111100001110001011011001,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000011010111,
    24'b111100011101111111010111,
    24'b111011001101101111010100,
    24'b111100001110010111011001,
    24'b010100000100100001001001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001000000101101010101010,
    24'b000000100110010111001010,
    24'b000000000110011111001010,
    24'b000000000110011111001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000100110100011001101,
    24'b000000110110011011001011,
    24'b000000100110010111010001,
    24'b000111100101100110100011,
    24'b000000000000110000101011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111011111110000111011001,
    24'b111100011110000111011010,
    24'b111100011110001011011010,
    24'b111100001110001011011001,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000111010110,
    24'b111100101110000111011000,
    24'b111011101101110011010100,
    24'b111100101110000111011010,
    24'b111011111110001111011010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001000100101101,
    24'b000111010101110110101101,
    24'b000000110110010011001100,
    24'b000000000110011011001110,
    24'b000000010110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000100110011111001111,
    24'b000000110110011011001100,
    24'b000001000110010011010010,
    24'b000110110101111110110001,
    24'b000000010001100000111111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111010111101111011010101,
    24'b111011111110000011011010,
    24'b111100001110000111011010,
    24'b111100001110001011011001,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100001101111111010111,
    24'b111100011110000111011010,
    24'b110111101101010011001101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001110001000101,
    24'b000101010101110110101111,
    24'b000000110110010111001101,
    24'b000000010110011011010010,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100011001110,
    24'b000000000110011111001110,
    24'b000000010110011111001111,
    24'b000000110110011011001110,
    24'b000000110110010011001110,
    24'b000101000110001010110111,
    24'b000010100010110101011011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110001001011101010110000,
    24'b111011111110001011011010,
    24'b111100001110001011011001,
    24'b111100001110001011011001,
    24'b111100011110000011011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110001011011000,
    24'b111100011110000011010111,
    24'b111100001101111111010111,
    24'b111101011110010011011101,
    24'b101101001010101110100101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000100000011100101110001,
    24'b000100100110010110111100,
    24'b000001000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110100011001110,
    24'b000000000110011111001110,
    24'b000000010110011011010000,
    24'b000000100110010011001111,
    24'b000000110110100011001111,
    24'b000011100110011011000000,
    24'b000011100100010110000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b011010100110000101011001,
    24'b111011111110010111011011,
    24'b111100011110010011011011,
    24'b111011101110000011010111,
    24'b111100111110001011011010,
    24'b111100011110000011010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111101111110010111011101,
    24'b111011011101110011010101,
    24'b010010110100010000111111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000110010101000010011010,
    24'b000001110110000111000000,
    24'b000000000110010111001111,
    24'b000000010110010111010001,
    24'b000000010110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110100011001100,
    24'b000000000110011011001100,
    24'b000000010110011011010000,
    24'b000000100110010011001111,
    24'b000001010110101011010011,
    24'b000010000110011111001001,
    24'b000110110101110110100011,
    24'b000000000000110100101101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111010101110001011011011,
    24'b111010111101111011010101,
    24'b111100111110010111011100,
    24'b111100001101111111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111010111101101011010010,
    24'b111110111110101011100011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000110100110111,
    24'b000111110101110010111000,
    24'b000000110110010111001100,
    24'b000000000110011011010010,
    24'b000000010110011111001101,
    24'b000000000110100011001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110100011001101,
    24'b000000000110011011001110,
    24'b000000010110011111010000,
    24'b000000100110010111010001,
    24'b000001100110101011010001,
    24'b000000010110010011001101,
    24'b000110110110011010111100,
    24'b000001000001111001001101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101111011011011010110001,
    24'b111100001110001111011011,
    24'b111100001110001011011001,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000011011000,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111011111110001011011001,
    24'b111100011110000111011001,
    24'b111100111110000011011001,
    24'b111101001110000111010111,
    24'b111100101110000111010110,
    24'b111101111110011111011110,
    24'b101111101010111110101011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000011100010100001011111,
    24'b000110010101111111000100,
    24'b000001010110101011010101,
    24'b000000100110100011010110,
    24'b000000010110100011001110,
    24'b000000000110011111001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000100110011111010001,
    24'b000001100110100011001101,
    24'b000000010110011111010101,
    24'b000100000110010111001011,
    24'b000100110100000010000001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b011000010101100001010111,
    24'b111010101101110111010110,
    24'b111100001110001011011001,
    24'b111011111101111011010101,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111011000,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000111010111,
    24'b111011101110001111010110,
    24'b111100011110001011011000,
    24'b111101001110000011011001,
    24'b111101001110000011010110,
    24'b111100001110001011010110,
    24'b111011101110010011011011,
    24'b001011000010001100100001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000101100100100110010000,
    24'b000011000101110111000110,
    24'b000001010110100111010110,
    24'b000000000110010111010101,
    24'b000000110110011111010001,
    24'b000000010110011011001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011111010000,
    24'b000000110110100011010010,
    24'b000000000110100011010010,
    24'b000000110110100011010110,
    24'b000010110110010111001011,
    24'b001000010101111110101011,
    24'b000000000001010000111000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111000001101011011001111,
    24'b111011001101111011010101,
    24'b111101001110001111011001,
    24'b111100111110001111010111,
    24'b111100111110000111010101,
    24'b111100101110001011010101,
    24'b111100101110000111010111,
    24'b111100011110001011010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110001011010100,
    24'b111100111110001011010011,
    24'b111100111110000011010011,
    24'b111100011110000011010111,
    24'b111011101110010011011110,
    24'b110100011100101111000110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001110001000100,
    24'b000111000110010010110100,
    24'b000001110110000111000100,
    24'b000001000110011011001111,
    24'b000000000110011011010100,
    24'b000000010110011011010001,
    24'b000000010110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000100110011111010001,
    24'b000000100110011111010001,
    24'b000001000110100111010011,
    24'b000000000110011011010100,
    24'b000000110110010011010000,
    24'b000010100110010011001011,
    24'b000101100110010110111100,
    24'b000001100011010001101011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b011110100111000001101010,
    24'b111100001110001111011011,
    24'b111100011110001111011001,
    24'b111100101110001011010101,
    24'b111100101110001011010011,
    24'b111100101110001011010101,
    24'b111100001110001011010101,
    24'b111100001110001011010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111101001110000011010111,
    24'b111100111110001011010010,
    24'b111100011110000111010001,
    24'b111100001110001011011000,
    24'b111011001110001011100001,
    24'b010100000100100101001001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000010100011111101111110,
    24'b000010010110011111000011,
    24'b000001000110011111000100,
    24'b000000110110010111001010,
    24'b000000000110100011010001,
    24'b000000010110010111010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110100011010111,
    24'b000010010110011111010000,
    24'b000010010110010111001001,
    24'b000010000110001011000001,
    24'b000110010101100110011110,
    24'b000000000001000000101100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111010011101111111011011,
    24'b111011111110001111011010,
    24'b111100011110001111010111,
    24'b111100011110000111010010,
    24'b111100101110001011010101,
    24'b111100011110001111010110,
    24'b111011111110000011010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000011011000,
    24'b111100111101111111011010,
    24'b111101101110010111011011,
    24'b111011011110000011010011,
    24'b111100001110000111011010,
    24'b110011111011111111000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001000100101010,
    24'b000101110101110110101101,
    24'b000000010110100011001110,
    24'b000000010110100011000110,
    24'b000000110110010111001000,
    24'b000000000110101011001111,
    24'b000000010110011111010010,
    24'b000000100110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000110110011011010101,
    24'b000001110110011011001111,
    24'b000001010110010011001001,
    24'b000010000110011111001100,
    24'b000101010110001010111000,
    24'b000001000010101001011110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b011011000110010001100010,
    24'b111010001101111011011000,
    24'b111011001110000011010101,
    24'b111011111110000111010100,
    24'b111100101110001011010101,
    24'b111100011110000011010110,
    24'b111100111110001011011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000011011001,
    24'b111100101110001111011011,
    24'b111011011110000011010111,
    24'b111100101110001011011100,
    24'b010101100100011001000110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000010110011100001101101,
    24'b000100100110001110111111,
    24'b000000000110101011010111,
    24'b000000010110100011001101,
    24'b000001000110011011001010,
    24'b000000000110100011001110,
    24'b000000000110011011010001,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000001010110011111010110,
    24'b000000110110011111010101,
    24'b000000010110011011001110,
    24'b000001100110011111001110,
    24'b000011000110010111001001,
    24'b000111000101101010100101,
    24'b000000000001001000110110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110010101100000110111101,
    24'b111011001110000111010111,
    24'b111011111110000111010101,
    24'b111100011110000011010110,
    24'b111101001110000111011010,
    24'b111100101101111111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010110,
    24'b111100111110000111010001,
    24'b111100001110001011011001,
    24'b111100101110010011100000,
    24'b110000011011001010101100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001011000111111,
    24'b000111100110000110110010,
    24'b000010110110010011000100,
    24'b000000100110010011010011,
    24'b000000000110010111010011,
    24'b000000100110011011001011,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110010011010101,
    24'b000000000110011011011000,
    24'b000000110110101011011000,
    24'b000000100110011111010000,
    24'b000001010110011011010000,
    24'b000101100110010110111110,
    24'b000011100011011001101111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001100000010100100101010,
    24'b111011011110001111011011,
    24'b111100001110000011010110,
    24'b111101001110001011011010,
    24'b111100101101111111011000,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010101,
    24'b111101001110001011001101,
    24'b111101001110011011011001,
    24'b111001101101101111010111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000110000101000,
    24'b000100010100000110000000,
    24'b000100010110010011000111,
    24'b000001100110001111000110,
    24'b000001000110001111010010,
    24'b000000110110011011011000,
    24'b000000010110100011001101,
    24'b000000010110011011001111,
    24'b000000000110011011010000,
    24'b000000000110011111001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010100,
    24'b000000100110010111010101,
    24'b000000100110010111010101,
    24'b000000000110100011010101,
    24'b000000000110101011001101,
    24'b000010010110010111000001,
    24'b000110000101110110110100,
    24'b000000000001011101000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b011110100110111101101100,
    24'b111101001110010111011110,
    24'b111011101110000011011010,
    24'b111110011110101111011110,
    24'b111101011110010111010011,
    24'b111101001110000111010110,
    24'b111100011110001011011001,
    24'b111100001110001011011001,
    24'b111100111110000111010101,
    24'b111101001110000011010100,
    24'b111100111110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110000111010110,
    24'b111011111110000111010100,
    24'b111101001110010011010111,
    24'b111100101110000111010100,
    24'b111100111110000111010010,
    24'b111100101110011011010101,
    24'b010110010101011101001100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001110101010001,
    24'b000110110110001010110110,
    24'b000001010110011011001101,
    24'b000000110110100011010010,
    24'b000000010110010111010000,
    24'b000000110110100011010010,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100011001110,
    24'b000000100110010111010000,
    24'b000000110110010111010011,
    24'b000000000110011011010100,
    24'b000000000110011111001110,
    24'b000010000110011011001010,
    24'b000100110110000011000001,
    24'b000110000100101110001110,
    24'b000000000000110000101101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101100111011000110101010,
    24'b111010111110101011011100,
    24'b111100101110000011010111,
    24'b111110001101111011011001,
    24'b111100101110000011010101,
    24'b111100011110001011011000,
    24'b111100011110000011010110,
    24'b111100111110000111010101,
    24'b111100111110000111010101,
    24'b111100111110000111010111,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110001011011000,
    24'b111100101110001011010110,
    24'b111100001110000011010100,
    24'b111011111101111011010011,
    24'b111100101110001111011111,
    24'b100111011001100010010110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000111100110011,
    24'b000101110101001010011010,
    24'b000011100110100111001000,
    24'b000000100110010111001110,
    24'b000001010110101011010100,
    24'b000000010110010111010000,
    24'b000000110110100011010010,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100011001100,
    24'b000000010110011011001110,
    24'b000001000110010011010010,
    24'b000000010110010111010100,
    24'b000000110110100111010101,
    24'b000001000110011111001111,
    24'b000011010110011011001101,
    24'b000101100110001010111111,
    24'b000011010011110101110111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110100011101001111001010,
    24'b111100101101111111011001,
    24'b111101101101110011010110,
    24'b111100011110000111011000,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111011000,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110001011010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111101001110001111011010,
    24'b111100111110001011011000,
    24'b111100111110000111010111,
    24'b111100111110001011011000,
    24'b111011111101111011010101,
    24'b111100111110010011011011,
    24'b110000111011100010110101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000101100100000101111101,
    24'b000011110110001110111110,
    24'b000000010110011111001111,
    24'b000000010110011111010001,
    24'b000000100110011111010001,
    24'b000000010110011011010000,
    24'b000000100110011111010001,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010001,
    24'b000000010110011011010001,
    24'b000000110110010111010011,
    24'b000000110110010111010100,
    24'b000000010110010111010001,
    24'b000000010110011111001110,
    24'b000001110110100111001110,
    24'b000010000110011111001100,
    24'b000101100101111110110001,
    24'b000010100010100001010001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001011010010010000100101,
    24'b111011011110001011011101,
    24'b111100101110001111011010,
    24'b111100101110010011011100,
    24'b111100101110000111010111,
    24'b111101001110000011010110,
    24'b111100101110000111011001,
    24'b111100001110001011011001,
    24'b111100011110000111010111,
    24'b111100101110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000111010110,
    24'b111100011110000111010110,
    24'b111100101110000111010111,
    24'b111100111110001011011000,
    24'b111100101110000011010110,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111011111101111011010110,
    24'b111011111110000011011001,
    24'b110110011100110011000101,
    24'b001010100010010000011001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000001100010101101100000,
    24'b000110010110000010110001,
    24'b000001110110010011001001,
    24'b000000000110100011010100,
    24'b000000010110011111010010,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010100,
    24'b000000000110011011010101,
    24'b000000000110011011010100,
    24'b000000010110011011010010,
    24'b000000010110011011010000,
    24'b000000010110011011001011,
    24'b000001000110011111001100,
    24'b000001000110101111000110,
    24'b000011010110011111000110,
    24'b000110100101010010101010,
    24'b000001000001101001000111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001010110010011100100110,
    24'b111000011110000011011011,
    24'b111011011110000011011010,
    24'b111101001101111111010101,
    24'b111110011110010011011001,
    24'b111100011110000011011001,
    24'b111011011110000111011011,
    24'b111011111110000111010111,
    24'b111100101110000011010010,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111101011110001111010111,
    24'b111011011101101111010000,
    24'b111101101110010011011000,
    24'b111100001101111111010101,
    24'b111001111101100011010001,
    24'b111001001101101111010110,
    24'b001011100010011100100100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001111001000111,
    24'b000101110110000110110010,
    24'b000010110110100011001000,
    24'b000001010110010111001010,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110100011010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000110110011011001110,
    24'b000001000110010111001110,
    24'b000001010110011111001000,
    24'b000001100110100011001111,
    24'b000011110110010111010001,
    24'b000101110100111110011111,
    24'b000000010001000100110011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001101100011011000111001,
    24'b111000101101011111010011,
    24'b111011111101101011010000,
    24'b111101001101110011010001,
    24'b111100001110000011011001,
    24'b111011001110000111011100,
    24'b111011111110000111010111,
    24'b111100101110000111010001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011101111111010001,
    24'b111101011110001111010101,
    24'b111100001101111011010001,
    24'b111101101110010111011100,
    24'b111000001101010111010000,
    24'b001010110010011000100110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000100001110001000010,
    24'b000110010101100010100001,
    24'b000010000110011011000110,
    24'b000000000110100011001110,
    24'b000000010110100011001101,
    24'b000000100110010111001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000000110011111001101,
    24'b000000000110100111001101,
    24'b000000000110100111001110,
    24'b000000010110011011001111,
    24'b000001010110010111010011,
    24'b000001100110001111010100,
    24'b000001010110001011010010,
    24'b000000110110010111010000,
    24'b000001000110101111010011,
    24'b000011010110001011000001,
    24'b000101110100110010001101,
    24'b000000010001010000101110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001111000011001000101110,
    24'b110110111100011110111101,
    24'b111100111101110111010100,
    24'b111100011110000111011100,
    24'b111011011110001111011110,
    24'b111100001110001011011000,
    24'b111100111110001011010010,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000111010111,
    24'b111100101110000111010110,
    24'b111100101110000111010110,
    24'b111100111110001011011000,
    24'b111011111101111111010110,
    24'b111011111101111111010110,
    24'b111100111110001011010111,
    24'b111101011110001111010100,
    24'b111100001101111111001111,
    24'b111101011110011011011001,
    24'b110010001011101010110011,
    24'b001011110010100100100101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001101001000010,
    24'b000110110101011010011101,
    24'b000011100110001011000001,
    24'b000001000110010111001001,
    24'b000000100110101111010010,
    24'b000000000110100011010001,
    24'b000000100110100011001111,
    24'b000000010110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010010,
    24'b000000100110011111010101,
    24'b000000010110011011010101,
    24'b000000100110011011010000,
    24'b000000110110010111001100,
    24'b000001000110010111001100,
    24'b000001100110010111001101,
    24'b000011100110001011000001,
    24'b000101010100111110010101,
    24'b000000000001010000111100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101110101011001110110001,
    24'b111010111101111011010111,
    24'b111100111110000111010111,
    24'b111101101110001111010110,
    24'b111101001110000111010011,
    24'b111100111110000111010101,
    24'b111100011110000111010111,
    24'b111100001110001011011001,
    24'b111100001110001011010110,
    24'b111100101110001011010100,
    24'b111100111110000111010101,
    24'b111101001110000111011001,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100111110000011011001,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100111110000111010101,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100011110001011011001,
    24'b111011101110000111010111,
    24'b111100111110001111010100,
    24'b111100011110000111010001,
    24'b111100101110001011011010,
    24'b111011101110000011011101,
    24'b111100001110000111011110,
    24'b111011111101111011011000,
    24'b111101001110000011011010,
    24'b111011101110010011010100,
    24'b101010001010000110011011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001101100111110,
    24'b000010000101010110100010,
    24'b000011100110010110111110,
    24'b000001100110010111000110,
    24'b000000010110011011001100,
    24'b000000000110011011001110,
    24'b000000000110100011001111,
    24'b000000000110011011001011,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110100011010010,
    24'b000000110110100011010010,
    24'b000001000110010111001101,
    24'b000000110110010011001101,
    24'b000001000110011011010001,
    24'b000001110110011111010000,
    24'b000100110110000010111010,
    24'b001000000101010010011001,
    24'b000000000001011001000010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100010111000001001111111,
    24'b111010011110000011011100,
    24'b111011111110001011011101,
    24'b111100011110000011010110,
    24'b111100011101111111010011,
    24'b111100111110001011011000,
    24'b111100001110000011010111,
    24'b111011111110000111010101,
    24'b111100101110001011010101,
    24'b111100111110000111010101,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010101,
    24'b111100111110000111010101,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111101001101111111011001,
    24'b111110001101111011011010,
    24'b111101111101111111010100,
    24'b111101011110000011010011,
    24'b111100101110000111010101,
    24'b111100111110001011011000,
    24'b111101101110010011010111,
    24'b111011101101101111001100,
    24'b111011001101101011010100,
    24'b011100110111000001100111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001101001000000,
    24'b000101010101100010011101,
    24'b000011000110010011000000,
    24'b000001110110010111000110,
    24'b000000110110011111001101,
    24'b000000010110011111010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110100011001111,
    24'b000000100110100111010100,
    24'b000000110110100011010100,
    24'b000000100110011011001110,
    24'b000000000110010111001111,
    24'b000000010110011011010010,
    24'b000010000110100111010001,
    24'b000011110110001011000010,
    24'b000110110101100110100111,
    24'b000000010010010001010011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010000110011111100111111,
    24'b110011101100011011000010,
    24'b111110011110101111100010,
    24'b111100011110000011011000,
    24'b111100011110000011010110,
    24'b111100101110000111010111,
    24'b111100101110001011010110,
    24'b111100101110001011010101,
    24'b111100101110000011010110,
    24'b111100111110000111010111,
    24'b111100011110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000111011001,
    24'b111100001110001011011000,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111011000,
    24'b111100111110000111011000,
    24'b111100111110000011010111,
    24'b111101111110000011011000,
    24'b111100101101110111011001,
    24'b111100001101110111010111,
    24'b111100011110011011011101,
    24'b110010111011111010110101,
    24'b010000000011000100101111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000001010010001101001100,
    24'b000110100101110110100011,
    24'b000010000110100111001010,
    24'b000001100110011111001101,
    24'b000001100110100011010000,
    24'b000000000110010111010001,
    24'b000000000110011011010100,
    24'b000000100110101011011001,
    24'b000000000110011011010101,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110100011001110,
    24'b000000000110011111001011,
    24'b000000000110011111010010,
    24'b000000010110100011010101,
    24'b000000100110011111001111,
    24'b000000000110011111001101,
    24'b000000000110011111001111,
    24'b000000000110011111010010,
    24'b000001000110010111010000,
    24'b000011000110010111000111,
    24'b000101100101110010101001,
    24'b000010010011010001101000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100001110111101101110011,
    24'b110111101101001011001111,
    24'b111100001110001111011011,
    24'b111011111101111111010101,
    24'b111100111110001111011001,
    24'b111101001110001111011011,
    24'b111100011110000111011000,
    24'b111100101110001111010110,
    24'b111100101110000011010110,
    24'b111100101110000011010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000011010111,
    24'b111100111110000111010111,
    24'b111101001110000011010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000111010111,
    24'b111100001110001011010111,
    24'b111100011110001011011001,
    24'b111100001110000111011001,
    24'b111100001110001011011001,
    24'b111100001110001011011001,
    24'b111100001110001011011000,
    24'b111100111110000111011000,
    24'b111100101101111111010110,
    24'b111100101110001111011000,
    24'b111010101110010111010101,
    24'b111010011110001011010110,
    24'b111100001110001111011011,
    24'b111100101110001011100000,
    24'b111000011101001011010011,
    24'b011100100110101001101100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000110100110000,
    24'b000010000011101101110101,
    24'b000110000110010010110011,
    24'b000001110110010011000011,
    24'b000000100110011111001111,
    24'b000000010110011111010001,
    24'b000000000110011011010010,
    24'b000000000110011011010011,
    24'b000000000110011111010100,
    24'b000000010110100111010110,
    24'b000000000110011011010011,
    24'b000000010110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000000110011111001101,
    24'b000000000110100011010001,
    24'b000000000110100011010010,
    24'b000000000110011111001110,
    24'b000000000110100011001011,
    24'b000000010110100011001010,
    24'b000000100110011011001100,
    24'b000000100110011011001111,
    24'b000000100110011011001101,
    24'b000001100110011011000110,
    24'b000101110110010110110110,
    24'b000101010100100010000000,
    24'b000000100001011100110101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100011001000010010000010,
    24'b111000111101100011010001,
    24'b111011111110000011011011,
    24'b111011111101111011011011,
    24'b111100101110010011011101,
    24'b111011101110000111010101,
    24'b111101111110001111011010,
    24'b111101011110000111011000,
    24'b111101001110000011010111,
    24'b111101001110000011010111,
    24'b111101001110000011010111,
    24'b111101001110000011010111,
    24'b111100111101111111010110,
    24'b111100111110000111011000,
    24'b111100111110000111011000,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100011110000011010111,
    24'b111100101110010011011010,
    24'b111011111110001011011001,
    24'b111011111110000111011000,
    24'b111100111110001111011010,
    24'b111011101101110111010100,
    24'b111101001101111111011001,
    24'b111100101110000111011011,
    24'b111011011110011011011101,
    24'b110100101101001011000101,
    24'b100000100111110101110000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001111101001100,
    24'b000011010101000010010111,
    24'b000010100110010110111100,
    24'b000001010110100011001100,
    24'b000000000110010111001110,
    24'b000000100110011011001110,
    24'b000000000110011111010000,
    24'b000000000110011111010001,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000110110011011001100,
    24'b000000110110011011001011,
    24'b000000010110011111001100,
    24'b000000000110011111001110,
    24'b000000000110010111001110,
    24'b000000110110001111000110,
    24'b000100100110001010111001,
    24'b001000010101110110100010,
    24'b000010100011000001100011,
    24'b000000000000111000110100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b011101110110101101101010,
    24'b110110011100110011001101,
    24'b111011101110001111100000,
    24'b111010111110001011010110,
    24'b111101011110010111011011,
    24'b111100101110000011010110,
    24'b111100001101111111010101,
    24'b111100101110000011010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100001110001011011001,
    24'b111100001110001011011001,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010110,
    24'b111100101110000111010101,
    24'b111100111110000011010101,
    24'b111101001110001011010110,
    24'b111011101110000011010101,
    24'b111011101110001011011001,
    24'b111011001110000111010111,
    24'b111100001110001111011011,
    24'b111011011101110111010111,
    24'b111110101110001011100010,
    24'b110100001011011110111011,
    24'b011011010110001101100001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010000111000101010,
    24'b000010110011011101100101,
    24'b000110000101110010101011,
    24'b000010110110100011001010,
    24'b000000110110101011001100,
    24'b000000100110100111001101,
    24'b000000010110011011010000,
    24'b000000010110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001101,
    24'b000000000110011111001101,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010100,
    24'b000000000110011011010100,
    24'b000000100110011011001111,
    24'b000000010110011011001110,
    24'b000000000110011011010100,
    24'b000000000110011011010101,
    24'b000000010110010111010011,
    24'b000000010110011011001110,
    24'b000000000110100011001110,
    24'b000000000110100011010000,
    24'b000000110110011011010000,
    24'b000001110110011111010000,
    24'b000001000110010111001111,
    24'b000000110110001011001110,
    24'b000101110110011011000111,
    24'b000110100101000110011100,
    24'b000001010010010101011010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001110110011000100101111,
    24'b100011101000011101111011,
    24'b111000101101100011001100,
    24'b111100011110011011011010,
    24'b111100001110011011011010,
    24'b111010001101110111010001,
    24'b111011101110001011010110,
    24'b111011111110010011011000,
    24'b111011111110001111010111,
    24'b111011111110001011011001,
    24'b111100001110001011011001,
    24'b111100001110001011011001,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111101001110000011010110,
    24'b111101001110000011010101,
    24'b111101011101111111010011,
    24'b111100111101111111010100,
    24'b111100101110000111010111,
    24'b111011001110000011010111,
    24'b111011101110010011011011,
    24'b110111001101000011001010,
    24'b100001100111100001110100,
    24'b001101110010101000101001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000110010101001011110,
    24'b000101110101110110100001,
    24'b000010110110011110111111,
    24'b000010100110000111001000,
    24'b000011010110011011001010,
    24'b000001100110011111000011,
    24'b000000100110100011001100,
    24'b000000000110011011010100,
    24'b000000000110011111010000,
    24'b000000000110011011010011,
    24'b000000010110011011010010,
    24'b000000010110011011010000,
    24'b000000010110011011001110,
    24'b000000000110011111001111,
    24'b000000000110011011010001,
    24'b000000000110011111010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010000,
    24'b000000100110100111010010,
    24'b000000100110100111010010,
    24'b000000010110011111010000,
    24'b000000100110011011001110,
    24'b000000110110010111001111,
    24'b000000110110010111010010,
    24'b000000100110001111010001,
    24'b000001110110011111001111,
    24'b000011110110100011001001,
    24'b000101110110001110111101,
    24'b000111010100011110011100,
    24'b000000110010000101011101,
    24'b000000010000111100101111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001010010010100100101010,
    24'b010111010101110001011001,
    24'b100100101000110010000111,
    24'b110001111100000010111011,
    24'b110101001100111011001001,
    24'b110111101101101111010100,
    24'b110111111101011011010000,
    24'b111010101101111011011000,
    24'b111010111101111011011100,
    24'b111011001101111111011100,
    24'b111011001101111111011100,
    24'b111001001101101011010101,
    24'b110111111101011011001111,
    24'b110101101100110111000010,
    24'b110010101100000110110111,
    24'b100100011000100110000000,
    24'b010101010100111101001001,
    24'b001010010010010100100010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001000000111011,
    24'b000001000010101001101011,
    24'b000110010101010010100100,
    24'b000100110101111010111000,
    24'b000010100110001011000011,
    24'b000000100110010111001011,
    24'b000001000110010111001111,
    24'b000001010110010011001111,
    24'b000000110110011011001111,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011001111,
    24'b000000010110100011010001,
    24'b000000010110100011010001,
    24'b000000000110011111001110,
    24'b000000000110011111001101,
    24'b000000010110011011001111,
    24'b000000010110011011010010,
    24'b000001000110011011010001,
    24'b000001000110010111001110,
    24'b000001000110011011001010,
    24'b000001100110100011001010,
    24'b000010110110101011000111,
    24'b000110000110011010111100,
    24'b000110100101001010011001,
    24'b000100000011001101101010,
    24'b000001100001011100111111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001011100010101100101011,
    24'b001011110010110100101100,
    24'b001011100010110100101100,
    24'b001011000010110100101011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000100010000001001000,
    24'b000011000011101101110010,
    24'b000101110101010010011110,
    24'b000100110101111110111000,
    24'b000011000110001111000110,
    24'b000000110110001111001001,
    24'b000000010110010011001001,
    24'b000000110110010111001100,
    24'b000001010110011111010001,
    24'b000001010110100011010110,
    24'b000001000110011111010110,
    24'b000000010110011111010011,
    24'b000000000110011111001111,
    24'b000000000110011111001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001101,
    24'b000000000110011111001111,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000110110011011010001,
    24'b000000110110011011001111,
    24'b000000010110011111001100,
    24'b000000000110111011001110,
    24'b000000110110100111001101,
    24'b000011100110011011001011,
    24'b000110000110000111000000,
    24'b000111110101101110101101,
    24'b000110010100111110001110,
    24'b000010010011100001101001,
    24'b000001110010000101000110,
    24'b000000000001000100110010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000101000101000,
    24'b000000000001010000111000,
    24'b000001000010010001010001,
    24'b000010100011001101101011,
    24'b000101010100111110010111,
    24'b000100010110000010111000,
    24'b000100010110011011000010,
    24'b000011000110100111001010,
    24'b000001000110011111001010,
    24'b000000000110010011001001,
    24'b000000000110100011001101,
    24'b000000000110011011001100,
    24'b000000110110011011001110,
    24'b000000110110010111010000,
    24'b000000110110011011010100,
    24'b000000110110011111010110,
    24'b000000010110011111010011,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011001111,
    24'b000000000110011011001111,
    24'b000000000110011111001111,
    24'b000000000110100011001101,
    24'b000000000110011111001111,
    24'b000000000110011011010010,
    24'b000000000110011011010100,
    24'b000000000110010111010001,
    24'b000000010110010111010001,
    24'b000000100110011111010001,
    24'b000000100110011111010000,
    24'b000000100110100111010000,
    24'b000000110110100111001111,
    24'b000000110110100011001101,
    24'b000000100110011011001011,
    24'b000001010110010011001001,
    24'b000010010110011011001000,
    24'b000100100110000110110110,
    24'b000101010101110110101011,
    24'b000101000101001010011001,
    24'b000011110100000001111100,
    24'b000100000011100001101010,
    24'b000000000010000001001100,
    24'b000000100001111101000101,
    24'b000000000001001000111101,
    24'b000000000000111100110110,
    24'b000000000000111000110001,
    24'b000000000001000000101111,
    24'b000000000000111100101111,
    24'b000000110001100100111100,
    24'b000001100001110101000101,
    24'b000010000010011101010111,
    24'b000001110010110101100111,
    24'b000100100011111101111111,
    24'b000101100101000010010110,
    24'b000101110101110110101000,
    24'b000100000110000110110100,
    24'b000010110110001011000000,
    24'b000010100110010111001100,
    24'b000001100110011011010000,
    24'b000000100110010011001100,
    24'b000000110110100011001101,
    24'b000000100110100011001100,
    24'b000000100110100011001100,
    24'b000000100110011011001010,
    24'b000000010110010111001010,
    24'b000000110110011011001110,
    24'b000000010110010011001111,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110100011001110,
    24'b000000000110011111001111,
    24'b000000000110011011010010,
    24'b000000000110011011010100,
    24'b000000000110011011010100,
    24'b000000000110011011010100,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110100011001110,
    24'b000000000110100111001100,
    24'b000000000110100111001011,
    24'b000000000110011111001111,
    24'b000000010110010111010101,
    24'b000000100110010011011000,
    24'b000000000110011011010000,
    24'b000000000110011011001011,
    24'b000001000110010111000110,
    24'b000010100110010010111111,
    24'b000011010110001110111000,
    24'b000100010110001110110101,
    24'b000101010110001110110010,
    24'b000110100110001110111000,
    24'b000110010110000110110010,
    24'b000110000101111110101101,
    24'b000110010101111110101011,
    24'b000110010101111110101011,
    24'b000101110110000010101111,
    24'b000110010110001010110101,
    24'b000100100110010010111110,
    24'b000011100110011011000111,
    24'b000010100110010011001000,
    24'b000001110110010011000111,
    24'b000001000110011111000110,
    24'b000000110110011111001001,
    24'b000000010110011111001100,
    24'b000000010110011011010000,
    24'b000000100110011011001111,
    24'b000000100110011011001100,
    24'b000000010110011111001100,
    24'b000000010110011111001100,
    24'b000000010110011111001100,
    24'b000000110110011011001110,
    24'b000000110110010111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010001,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011011010010,
    24'b000000100110010111010011,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011111001011,
    24'b000000100110011111001000,
    24'b000000110110011011001010,
    24'b000000100110011111001010,
    24'b000000010110011011001010,
    24'b000000000110011011001100,
    24'b000000000110011111001110,
    24'b000000010110100011010000,
    24'b000000010110100011010000,
    24'b000001000110100111001101,
    24'b000001000110100011001001,
    24'b000001000110011111000111,
    24'b000001000110100011000110,
    24'b000001000110100011000110,
    24'b000001000110100111001001,
    24'b000000110110100011001001,
    24'b000000110110011011001000,
    24'b000001010110010011001011,
    24'b000001000110011111001111,
    24'b000000100110100011010010,
    24'b000000010110100111001111,
    24'b000000000110100111001111,
    24'b000000000110011111010001,
    24'b000000000110011011010010,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010011,
    24'b000000000110011111010100,
    24'b000000000110011011010101,
    24'b000000000110011011010101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011001111,
    24'b000000010110011111001111,
    24'b000000010110011111001111,
    24'b000000010110011111010000,
    24'b000000000110011011010001,
    24'b000000100110011011010001,
    24'b000000010110011011010011,
    24'b000000010110011011010011,
    24'b000000000110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111001111,
    24'b000000000110100011001101,
    24'b000000010110011111001111,
    24'b000000100110011111001111,
    24'b000000000110011011010000,
    24'b000000000110010111010000,
    24'b000000100110011111010001,
    24'b000000110110011011010001,
    24'b000001000110011011010000,
    24'b000000110110011111001100,
    24'b000000110110100011001110,
    24'b000001010110011111001111,
    24'b000001010110011111001111,
    24'b000001000110011011001110,
    24'b000000110110010111001100,
    24'b000000100110011111001100,
    24'b000000110110011111001111,
    24'b000000110110011011010000,
    24'b000000100110011111010100,
    24'b000000010110100011010100,
    24'b000000000110100011001111,
    24'b000000000110011111001110,
    24'b000000100110011011010000,
    24'b000000010110010111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010001,
    24'b000000010110011011010011,
    24'b000000010110011011010011,
    24'b000000010110011111010001,
    24'b000000010110011111001110,
    24'b000000010110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010010,
    24'b000000000110011111010011,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110010111010001,
    24'b000000100110011011010001,
    24'b000000100110011011010000,
    24'b000000110110010111010001,
    24'b000000110110010111010010,
    24'b000001000110010111010001,
    24'b000001000110010111010001,
    24'b000000110110010111010010,
    24'b000000110110010111010010,
    24'b000000100110011111010010,
    24'b000000010110011011010100,
    24'b000000000110011011010011,
    24'b000000000110011111010001,
    24'b000000000110011011001110,
    24'b000000000110011111001101,
    24'b000000000110011111001100,
    24'b000000100110011011001101,
    24'b000000010110010111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011001111,
    24'b000000010110011111001101,
    24'b000000000110011111001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010011,
    24'b000000010110011111010011,
    24'b000000010110011111010011,
    24'b000000100110011111010011,
    24'b000000100110011111010011,
    24'b000001000110011011010001,
    24'b000001000110011011010001,
    24'b000001000110011011010001,
    24'b000000010110011011010010,
    24'b000000000110011011010100,
    24'b000000010110011011010010,
    24'b000000010110011011010000,
    24'b000000010110011011001101,
    24'b000000010110011111001011,
    24'b000000000110100011001011,
    24'b000000000110011111001100,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000000110011011010010,
    24'b000000000110010111010001,
    24'b000000000110010111010001,
    24'b000000000110010111001111,
    24'b000000000110010111001111,
    24'b000000010110011011010000,
    24'b000000010110011111010100,
    24'b000000000110100011010101,
    24'b000000010110011111010100,
    24'b000000010110011011010000,
    24'b000000010110011011001110,
    24'b000000010110011111001100,
    24'b000000010110100011001101,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000000110011111001110,
    24'b000000000110011111001100,
    24'b000000000110011111001110,
    24'b000000100110100111010000,
    24'b000000100110100111010010,
    24'b000000000110100111010010,
    24'b000000000110100011010011,
    24'b000000000110100011010011,
    24'b000000010110100011010001,
    24'b000000010110100011010001,
    24'b000000010110100011010001,
    24'b000000000110100111010101,
    24'b000000000110100111010110,
    24'b000000010110011111010011,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110100011001111,
    24'b000000010110100011001111,
    24'b000000010110100011001111,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000
};

assign mem = memory;

endmodule
