module sprite_tile(output logic [23:0] mem [0:4899]);

logic [23:0] memory [0:4899] = '{
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011011010001,
    24'b000000010110011011010001,
    24'b000000010110011011010000,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011001111,
    24'b000000000110011011001111,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010001,
    24'b000000010110011011010001,
    24'b000000010110011011010001,
    24'b000000010110011011010001,
    24'b000000010110011011010001,
    24'b000000000110100011001110,
    24'b000000000110100011001110,
    24'b000000000110011111001110,
    24'b000000010110100011001101,
    24'b000000000110011111001110,
    24'b000000000110011111001101,
    24'b000000000110011111001100,
    24'b000000010110011111001100,
    24'b000000010110011111001100,
    24'b000000000110011111001100,
    24'b000000000110100011001100,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000100110011111001111,
    24'b000000100110011111001111,
    24'b000000100110011111010001,
    24'b000000010110011011010000,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000000110100011010011,
    24'b000000000110100011010011,
    24'b000000000110100011010001,
    24'b000000000110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000010110100011010001,
    24'b000000010110100011001111,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000010110011011001111,
    24'b000000010110011011001111,
    24'b000000100110011011001110,
    24'b000000010110011011001111,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111001110,
    24'b000000100110100011001110,
    24'b000000010110011011001111,
    24'b000000100110011111010010,
    24'b000000100110011011010100,
    24'b000000100110011011010101,
    24'b000000000110011111010011,
    24'b000000000110100011010010,
    24'b000000010110011111010001,
    24'b000000010110011111010000,
    24'b000000110110011111001111,
    24'b000000100110011111001111,
    24'b000000010110011111001111,
    24'b000000010110011111001100,
    24'b000000010110011111001100,
    24'b000000100110100111001110,
    24'b000000110110100111010010,
    24'b000001000110100111010100,
    24'b000000100110011111010010,
    24'b000000100110100011010100,
    24'b000000010110011111010011,
    24'b000000100110011111010100,
    24'b000000100110011111010100,
    24'b000000100110011111010011,
    24'b000001000110011011010011,
    24'b000001000110011011010011,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111001100,
    24'b000000000110011011001011,
    24'b000000010110011011001110,
    24'b000000010110011011010010,
    24'b000000010110010111010100,
    24'b000000000110010011010100,
    24'b000000010110100011010001,
    24'b000000010110011011001111,
    24'b000001000110011111001111,
    24'b000001000110011011001100,
    24'b000001000110010111001011,
    24'b000001000110010111001011,
    24'b000001010110011011001011,
    24'b000001000110010111000110,
    24'b000001000110010111000101,
    24'b000001010110011011001000,
    24'b000001010110010111001011,
    24'b000001000110010111001011,
    24'b000001000110011011001011,
    24'b000000110110011011001101,
    24'b000001000110011011010000,
    24'b000000110110010111010000,
    24'b000000010110011011010001,
    24'b000000110110011011010000,
    24'b000001000110011011010001,
    24'b000001000110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000100110011111010000,
    24'b000000010110011011001110,
    24'b000000000110010111001110,
    24'b000000010110011111010001,
    24'b000001000110101111010111,
    24'b000000110110100111010100,
    24'b000000100110010011001100,
    24'b000001000110011011001011,
    24'b000001110110011011000111,
    24'b000010110110001111000001,
    24'b000100100110001111000000,
    24'b000100110110001010111100,
    24'b000100000101111010110110,
    24'b000100010101101110110011,
    24'b000100000101101110101111,
    24'b000100000101101110101101,
    24'b000100000101101110101111,
    24'b000101000101111010110111,
    24'b000011110110010110111100,
    24'b000010010110001010111010,
    24'b000010010110010011000001,
    24'b000001100110010111000101,
    24'b000001000110010011001010,
    24'b000001010110010111001111,
    24'b000001000110011111001011,
    24'b000001000110011111001111,
    24'b000000110110100011010001,
    24'b000000010110011011001111,
    24'b000000000110011111001111,
    24'b000000000110100011010001,
    24'b000000000110011111010000,
    24'b000000100110011011001110,
    24'b000000000110100011010010,
    24'b000000000110100011010010,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110100011010010,
    24'b000000000110011111001111,
    24'b000000110110010111001010,
    24'b000000000110010111001111,
    24'b000000110110100111010001,
    24'b000001000110010011001001,
    24'b000011000110100011001011,
    24'b000001110110000111000100,
    24'b000100010110011011000110,
    24'b000101010110001110111011,
    24'b001000100101011110011100,
    24'b000100010011111001111000,
    24'b000001110010011101010110,
    24'b000000000001011100111010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001000000110011,
    24'b000000000001110101001001,
    24'b000010010011010101101000,
    24'b000101000100111110001100,
    24'b000101110101111010101001,
    24'b000100110110000110111010,
    24'b000011110110001111001001,
    24'b000001000110010111001100,
    24'b000000100110100111001111,
    24'b000001000110101011010000,
    24'b000000010110011011010000,
    24'b000000000110011011010100,
    24'b000000000110011111001111,
    24'b000000000110100011001011,
    24'b000000000110100011010001,
    24'b000000000110011011010010,
    24'b000000110110011011001100,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000000110011011010010,
    24'b000000110110011011001101,
    24'b000001010110011011001101,
    24'b000000000110100011010100,
    24'b000000000110100011010101,
    24'b000010110110010111001000,
    24'b000111110110000010110000,
    24'b001000000100110110001010,
    24'b000001110010010001010011,
    24'b000000010000111100110011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000100001001100110010,
    24'b000011010011100101111000,
    24'b000111010101101110110001,
    24'b000110000110100011001100,
    24'b000010100110010011001100,
    24'b000000110110011111001001,
    24'b000000100110011011001011,
    24'b000000110110011111001010,
    24'b000000100110011011001000,
    24'b000000100110010111001100,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111001101,
    24'b000001010110100011001110,
    24'b000000000110011011010111,
    24'b000000010110101011011111,
    24'b000011010110001111000111,
    24'b000111100101110110101110,
    24'b000011110011101001111001,
    24'b000000000001000000111000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001011010010010100100011,
    24'b011101100110101101100100,
    24'b101010101001110110010101,
    24'b110100001100001110111001,
    24'b110111101101000011001000,
    24'b111001001101010111001111,
    24'b111001101101011011010000,
    24'b111001101101011011010010,
    24'b111000101101001011001111,
    24'b110111011100110011001000,
    24'b101101101011000110100110,
    24'b100011001000100010000001,
    24'b010100010100110001001010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000001000010010001010110,
    24'b000101000100111110010111,
    24'b000011010110001010111110,
    24'b000001000110101011001100,
    24'b000000110110010111001010,
    24'b000000010110001011001100,
    24'b000000000110100011010011,
    24'b000000010110110011011000,
    24'b000000010110010111010100,
    24'b000000100110010111010000,
    24'b000000100110011011010001,
    24'b000000010110011011010000,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010000,
    24'b000000000110011111001111,
    24'b000000000110011111001100,
    24'b000010000110011111001000,
    24'b000010100110011011001010,
    24'b000100010110001110111101,
    24'b000011100011111001111101,
    24'b000000010001000100101101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010100110100101101001101,
    24'b101101111010111010110000,
    24'b111000111101011011010000,
    24'b111011101101111111011001,
    24'b111100011110001011011010,
    24'b111100011110001011011001,
    24'b111100101110001011011000,
    24'b111100011110001111011000,
    24'b111011111110000111010101,
    24'b111100001110001011010110,
    24'b111100001110001011010111,
    24'b111100001110001011011000,
    24'b111100011110001111011001,
    24'b111100001110000011010110,
    24'b111100001110000011011011,
    24'b111011011110000011011101,
    24'b111011001110010111011101,
    24'b110011111100110011000011,
    24'b011110010111100001110000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000001100010010001010101,
    24'b000101000101011110100010,
    24'b000010100110100111000100,
    24'b000000100110110011010100,
    24'b000001000110010011010010,
    24'b000010100110000111001010,
    24'b000001010110011011000110,
    24'b000000110110011011001110,
    24'b000000110110011011001110,
    24'b000000010110011011010000,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000010110100011010001,
    24'b000000010110011111010001,
    24'b000001010110010111010001,
    24'b000011100110010111001001,
    24'b000101110100111010010100,
    24'b000000100001010000110010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100010100111111101111010,
    24'b110111111101010111001100,
    24'b111011101110001111011100,
    24'b111100101110001111011011,
    24'b111011001101111111010101,
    24'b111100101110010011011011,
    24'b111100011110001011011001,
    24'b111101001110010011011011,
    24'b111100011110000011010110,
    24'b111011111101110111010010,
    24'b111100011110000111010001,
    24'b111100111110000111010110,
    24'b111100111110000111010111,
    24'b111100111110001011010111,
    24'b111100111110000111010101,
    24'b111100001110000111010110,
    24'b111011101101111111011010,
    24'b111100101110001111011110,
    24'b111011111110000111011000,
    24'b111011101110000111010011,
    24'b111100011110010011010111,
    24'b111100011110001011011010,
    24'b101110111011001110101111,
    24'b010000100011110100111100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000010100011010001101001,
    24'b000101110110000010110110,
    24'b000011000110011011001111,
    24'b000001000110010111010000,
    24'b000000010110100011010010,
    24'b000001000110010111001110,
    24'b000000110110010111001110,
    24'b000000110110010111010000,
    24'b000000100110011111010001,
    24'b000000000110011111010001,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011011001110,
    24'b000000010110011011001110,
    24'b000000000110010111001111,
    24'b000000000110011011010010,
    24'b000000000110011111010100,
    24'b000000010110011011001101,
    24'b000000000110011111010100,
    24'b000000000110100011010100,
    24'b000001100110100011001110,
    24'b000000110110100011010001,
    24'b000101100110001110110011,
    24'b000011100011001101101110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100001000111100001110110,
    24'b111011011101110111010101,
    24'b111101001110001111011010,
    24'b111100011110001011011000,
    24'b111100011110001011011000,
    24'b111100011110001011010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100111110000111010101,
    24'b111100101110000111010110,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100101110000111011000,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010110,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111101001110000111100001,
    24'b111101001110001111011011,
    24'b111100101110001111010110,
    24'b110001011011100110101111,
    24'b001100110010101000100111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000110001010100111011,
    24'b000110110101100010100011,
    24'b000010100110011011001011,
    24'b000001010110100011010000,
    24'b000000110110101111010100,
    24'b000000000110011011010001,
    24'b000000000110011111010010,
    24'b000001010110100011010000,
    24'b000000000110011011001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011011001110,
    24'b000000100110011111001111,
    24'b000000010110011011010000,
    24'b000000000110011011010011,
    24'b000000010110011111001101,
    24'b000000010110011011001110,
    24'b000000010110011111001100,
    24'b000000000110011111010000,
    24'b000001010110011011001001,
    24'b000110010101110010101000,
    24'b000000100010001101010100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001111010011101001000110,
    24'b111000011101011011010101,
    24'b111011011101110111010010,
    24'b111100001101111111010101,
    24'b111100111110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100011110000111011101,
    24'b111101101110001111011100,
    24'b111100011101111111010100,
    24'b111100011110001111011010,
    24'b111100001110010111011110,
    24'b100110011000111110001011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000101000101001,
    24'b000101000100010010000000,
    24'b000101010110011110111111,
    24'b000000000110101011010101,
    24'b000001010110010111001101,
    24'b000010000110010111001100,
    24'b000000110110100111001111,
    24'b000000000110011111010000,
    24'b000000010110011011001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001111,
    24'b000000010110011011010000,
    24'b000000100110011111010001,
    24'b000000110110011011001100,
    24'b000000000110011111010010,
    24'b000000010110011011001110,
    24'b000001010110000111000001,
    24'b000101000101011010011111,
    24'b000000100001011100111011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b100101111000100110000100,
    24'b111010011110001011010001,
    24'b111100111110010011011101,
    24'b111100101101111011011000,
    24'b111100101110000111010111,
    24'b111100001101111111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111011111110001011010101,
    24'b111100111110001011011010,
    24'b111101001110000111011010,
    24'b111110001110011111011111,
    24'b111011001101111011010001,
    24'b111011101101110011001101,
    24'b110111001101010111001101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000011000011100101110000,
    24'b000011010110010110111111,
    24'b000011000110001011001100,
    24'b000000110110001111010001,
    24'b000000000110101111010000,
    24'b000000000110011111001110,
    24'b000000100110010111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110010111010000,
    24'b000000100110011111010000,
    24'b000000010110011111010100,
    24'b000000010110011011010100,
    24'b000001100110010011001110,
    24'b001000110101101110100011,
    24'b000000000000110100101100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110010011100000010111001,
    24'b111100101110010111011110,
    24'b111100001110010111011110,
    24'b111101001110001011011000,
    24'b111100111110000111010100,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010100,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100001110000011010001,
    24'b111011011110010011011000,
    24'b111010111110100011100001,
    24'b010010000100010101000001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000100110011101101101110,
    24'b000100110110001111000001,
    24'b000000000110100111011011,
    24'b000000100110101111010011,
    24'b000000110110011011001101,
    24'b000000010110011111010010,
    24'b000000000110011111001110,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010001,
    24'b000000000110010111010001,
    24'b000000110110100011010010,
    24'b000001000110011011001110,
    24'b000000010110011011010000,
    24'b000010100110010111000101,
    24'b000111100101111010101011,
    24'b000000010001001000110110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110101101100111011000110,
    24'b111100011110010011011110,
    24'b111010101101110011010011,
    24'b111100101110010011011001,
    24'b111011111110000111010110,
    24'b111100101110000111010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010110,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110000111010110,
    24'b111100011110001111011001,
    24'b111100001110001011011001,
    24'b111010111101111111011000,
    24'b111010101110000111100000,
    24'b011010010110010001100101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000010100011110101110010,
    24'b000011100110011010111111,
    24'b000010000110010011001111,
    24'b000001010110010111010000,
    24'b000000000110011111010011,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010011,
    24'b000000110110011111001111,
    24'b000001010110011111001110,
    24'b000001010110011111001000,
    24'b000101110110001110110001,
    24'b000000000001001100111000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110101111101000011000011,
    24'b111101001110001111010101,
    24'b111100011101110111010011,
    24'b111101001101111111010010,
    24'b111100111110001011010001,
    24'b111100011110001011011000,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000011011001,
    24'b111100111110000111010110,
    24'b111100101110001011010011,
    24'b111100101110001011010101,
    24'b111100101110000111011001,
    24'b111100011110001011011010,
    24'b111101001110001111011011,
    24'b111110011110001111011100,
    24'b111101011101111011010110,
    24'b111100001110000011011010,
    24'b011011000110010101100010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000110100100111010000100,
    24'b000011110101111111000111,
    24'b000000100110010111010011,
    24'b000000000110011111010001,
    24'b000000010110011111010101,
    24'b000000000110011011010011,
    24'b000000000110011111010001,
    24'b000000000110011111001101,
    24'b000000000110011111001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010001,
    24'b000000010110011011001110,
    24'b000000010110011011001111,
    24'b000000000110011111010100,
    24'b000010000110100011001110,
    24'b000000110110010111001011,
    24'b000100000110010111000011,
    24'b000001100010100101011110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110100001100100010111111,
    24'b111100001110001111010101,
    24'b111100001110000011010001,
    24'b111100101110001011010101,
    24'b111100011110000111010100,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110000111010111,
    24'b111100101110000011010110,
    24'b111011111101110011010101,
    24'b111100001101110011010110,
    24'b001111010011010100111000,
    24'b000000000000000000000000,
    24'b000000000000111100101001,
    24'b000110110101100110100110,
    24'b000010000110101011001000,
    24'b000001110110011011010000,
    24'b000001000110100011010110,
    24'b000000000110011011011000,
    24'b000000000110011111010001,
    24'b000000010110100011001001,
    24'b000000000110011111010000,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110100011001011,
    24'b000000010110011011001111,
    24'b000000000110001111001101,
    24'b000010100110001110111011,
    24'b000100000100001101110111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101110101010110010100101,
    24'b111100111110011011100000,
    24'b111011101101110011010011,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110001011010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100011110000111010111,
    24'b111100101110000111010111,
    24'b111101111110011011011100,
    24'b111101011110010011011100,
    24'b111011001101110111010001,
    24'b001010110010010000100110,
    24'b000000000000000000000000,
    24'b000000000001100100111011,
    24'b000101110110000110111000,
    24'b000010110110011111001001,
    24'b000001000110001111010001,
    24'b000000110110011111010000,
    24'b000000110110010111010000,
    24'b000000100110010111010011,
    24'b000000000110011011010101,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000000110011111010010,
    24'b000000000110100011001101,
    24'b000001000110010011010001,
    24'b000001010110010011010010,
    24'b000101100101101110100011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b011000010101001101001011,
    24'b111100001110010011011011,
    24'b111011111110000111011001,
    24'b111100111110000111010101,
    24'b111100001110000011010011,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111011111110000111010110,
    24'b111011011101111111010100,
    24'b111100011110001011010111,
    24'b111100011110000011001110,
    24'b111000111101011011011010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000010000011010001101010,
    24'b000010010101111110111111,
    24'b000001100110100111010111,
    24'b000000010110011011001111,
    24'b000000110110010111010000,
    24'b000000110110010111010100,
    24'b000000000110011111010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010100,
    24'b000000010110010111010100,
    24'b000001010110010011010010,
    24'b000101000110001111000000,
    24'b000001110010101001011110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111100011110011011100000,
    24'b111010101110000011010111,
    24'b111100001110010011011001,
    24'b111100101110001011010100,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111011011101111011010000,
    24'b111011101110000011011011,
    24'b100011101000001110000010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000110000101101110101001,
    24'b000001010110100011001101,
    24'b000000000110011111010010,
    24'b000000010110100011010001,
    24'b000000110110011011001100,
    24'b000000010110011111001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100011001110,
    24'b000000110110011011001011,
    24'b000001010110001111010101,
    24'b000000110110010011001101,
    24'b000110010101011010010101,
    24'b000000000000110100101011,
    24'b000000000000000000000000,
    24'b110001111011111010111100,
    24'b111001111101110011010110,
    24'b111100001110001011011010,
    24'b111011111101111111010101,
    24'b111100111110000111011000,
    24'b111100101110000111011001,
    24'b111100101110000111011001,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000011011000,
    24'b111100111110000011011001,
    24'b111100111110000011011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100001110001011010111,
    24'b111101011110000111011000,
    24'b111010001110001111011001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000110010010101000110,
    24'b000101100110011110111011,
    24'b000001010110010111010101,
    24'b000000000110100011010010,
    24'b000000000110100011000111,
    24'b000000010110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001100,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111001101,
    24'b000000100110011111010010,
    24'b000000000110011111010011,
    24'b000001000110100011001010,
    24'b000000110110000111010000,
    24'b000011110110010111000010,
    24'b000001100010001001001001,
    24'b000000000000000000000000,
    24'b001110100011010000110010,
    24'b111100001110010111100000,
    24'b111100011110001011011011,
    24'b111100001110001011010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010110,
    24'b111100011110000011010110,
    24'b111100111110000111011010,
    24'b111011011110001111011010,
    24'b110001011011100110110111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001000010110001010100010,
    24'b000001100110000111001110,
    24'b000001100110011011001111,
    24'b000000000110101011010100,
    24'b000000000110011111010011,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001100,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001100,
    24'b000000100110011011010010,
    24'b000000100110010111010011,
    24'b000000100110101011000111,
    24'b000011110110110111010010,
    24'b000111110101101110100110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110011011100010010111110,
    24'b111100111110010111011101,
    24'b111100111110001011011001,
    24'b111100001110001011010101,
    24'b111100001110001011010101,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110001111010110,
    24'b111100011110001111011011,
    24'b111011111101111111011000,
    24'b111100001110001011011011,
    24'b001100000010101000100110,
    24'b000000000000000000000000,
    24'b000000010010001101010010,
    24'b000101110110101011001010,
    24'b000010010110001111001100,
    24'b000000010110011111010100,
    24'b000000000110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000010110011011010010,
    24'b000001000110010011010010,
    24'b000000000110101111000101,
    24'b000010010110001111000001,
    24'b000010110010100101011101,
    24'b000000000000000000000000,
    24'b001011000010100000101000,
    24'b111011011110001011011000,
    24'b111100011110000011010100,
    24'b111100011101111111010011,
    24'b111100001110001011010101,
    24'b111011111110001111010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111011101110000111011001,
    24'b111011101101111111011000,
    24'b111100001110000011011000,
    24'b101110111011001010101110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001000100110000110101101,
    24'b000010100110011011010000,
    24'b000001010110010011001111,
    24'b000000000110011011001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000001000110010111010000,
    24'b000000000110101111001010,
    24'b000101100110100010111001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101001011010001010100011,
    24'b111011011110001111010111,
    24'b111100101110000111010100,
    24'b111101001110000111010011,
    24'b111100011110001011010101,
    24'b111100001110001011010110,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100001110001011011001,
    24'b111100101110000111011001,
    24'b111100111110001011011001,
    24'b111011111110001111011101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000111000100101010000100,
    24'b000010000110010011001100,
    24'b000001000110010111010000,
    24'b000000000110011111010001,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111001110,
    24'b000000000110011111010001,
    24'b000000000110011011010100,
    24'b000000010110011011010000,
    24'b000000110110011011001100,
    24'b000000110110100011001111,
    24'b000110000101011110010111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111010101110001011011110,
    24'b111100011110010011011011,
    24'b111100101110000111010111,
    24'b111100111101111111010101,
    24'b111100101110000111010101,
    24'b111100101110000111010111,
    24'b111100111110000011011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010101,
    24'b111100011110000111011000,
    24'b111100101110000111010111,
    24'b111101001110001011010111,
    24'b111011001101111111010111,
    24'b011011110110100001100100,
    24'b000000000000000000000000,
    24'b000000000001010000111111,
    24'b000100100110010111000001,
    24'b000000110110011111010001,
    24'b000000000110011111010011,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111001100,
    24'b000000000110011111010001,
    24'b000000000110011011010110,
    24'b000000010110011011010000,
    24'b000000100110011111001000,
    24'b000011000110010011001111,
    24'b000000110010110101011010,
    24'b000000000000000000000000,
    24'b010001000100000101000001,
    24'b111101011110010011010111,
    24'b111100001110010011011101,
    24'b111100001110000111011001,
    24'b111101001110000011010111,
    24'b111100111110000111010111,
    24'b111100111110000011011000,
    24'b111101001110000011011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111011000,
    24'b111100111110000111010111,
    24'b111100111110000011010100,
    24'b111011101110000011011000,
    24'b110110101101000011001011,
    24'b000000000000000000000000,
    24'b000000000001000000101111,
    24'b000110010101111110101011,
    24'b000000110110011011001100,
    24'b000000100110011011001101,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011011010001,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000010110011011010000,
    24'b000000010110011011001110,
    24'b000011000110010010111101,
    24'b000000010001000100101100,
    24'b000000000000000000000000,
    24'b100110101001011110010101,
    24'b111101011110010011011001,
    24'b111100011110010111011010,
    24'b111011101110000111010101,
    24'b111101011110001111011001,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111011011101110011010100,
    24'b111011101110001011011011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000111010101011010010011,
    24'b000001110110100011001010,
    24'b000000100110011111010110,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110011011010001,
    24'b000000010110011011010000,
    24'b000000010110011011001110,
    24'b000100010101111110110001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110110001101000111001011,
    24'b111100001101111011010001,
    24'b111100111110010111011010,
    24'b111100001110001011010111,
    24'b111100001101111111010101,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000011011000,
    24'b111100001101111111010111,
    24'b111011111110000111011010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000011100011110101110100,
    24'b000010010110011111000110,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000110110011011001101,
    24'b000111110101111110100110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111011001110000011011000,
    24'b111101101110001111010110,
    24'b111011111101111111010101,
    24'b111100001110001011010111,
    24'b111100111110001011011000,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111011101101110111010101,
    24'b111100111110000111011001,
    24'b100000110111010001101110,
    24'b000000000000000000000000,
    24'b000000000001111001001100,
    24'b000010110110010010111111,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000010110011011001111,
    24'b000000100110011111010001,
    24'b000001010110010111001011,
    24'b001000100101001010001111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111100101110000111010111,
    24'b111101001110001011011000,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100011110001011010111,
    24'b111100011110001011010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100111110001011011010,
    24'b111100001101110111010011,
    24'b110100101100010010111110,
    24'b000000000000000000000000,
    24'b000000000000111100110011,
    24'b000011100110000110111100,
    24'b000000000110011111001110,
    24'b000000000110011111010001,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011011001111,
    24'b000000010110011011010010,
    24'b000001110110011011001101,
    24'b000110010011111101110011,
    24'b000000000000000000000000,
    24'b001010000010001000100001,
    24'b111100101110000011010101,
    24'b111100111110001011011011,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100001101111111010111,
    24'b111101011110001011011000,
    24'b110111111101010111001111,
    24'b000000000000000000000000,
    24'b000000000000101100101001,
    24'b000100100110001010111011,
    24'b000000000110011111001110,
    24'b000000000110011011010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111001111,
    24'b000000010110011111001111,
    24'b000000010110011011001111,
    24'b000010000110011111001100,
    24'b000011110011001001100101,
    24'b000000000000000000000000,
    24'b010100100100111001001100,
    24'b111100111110001111010110,
    24'b111011111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000011011000,
    24'b111100101110000111011001,
    24'b111100101110000111010110,
    24'b111000111101101011010010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000101010110001010111000,
    24'b000000100110011011010000,
    24'b000000010110011011010001,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010000,
    24'b000001010110011111010010,
    24'b000010010110011111001100,
    24'b000001100010110001011111,
    24'b000000000000000000000000,
    24'b011001100110001001011110,
    24'b111100101110001111010111,
    24'b111100101110001011010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011011000,
    24'b111001111101111111010110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000101000110001010110000,
    24'b000000100110010111010001,
    24'b000000010110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011111010000,
    24'b000001010110011111010100,
    24'b000010010110011111001101,
    24'b000001100010100101011100,
    24'b000000000000000000000000,
    24'b011010000110001101100000,
    24'b111101001110001011011000,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111011111110001111010111,
    24'b111001101110000011010110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000101110110000110110000,
    24'b000000000110011011001111,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110011011001110,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000100110100011010010,
    24'b000001000110011011010011,
    24'b000010010110011111001101,
    24'b000001110010110101011111,
    24'b000000000000000000000000,
    24'b010110110101010001010010,
    24'b111101001110000111011000,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100011110000011010110,
    24'b111100001110001011010111,
    24'b111100001110001111011000,
    24'b111001011101111111010100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000101000110000010110001,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000001010110011011010100,
    24'b000010000110011111001110,
    24'b000100010011101101101111,
    24'b000000000000000000000000,
    24'b001110010011001000110000,
    24'b111100101110000011010111,
    24'b111100011110000011010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111000011101101011010010,
    24'b000000000000000000000000,
    24'b000000000000100000101110,
    24'b000100100110000110110111,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011111010000,
    24'b000000010110011111010000,
    24'b000001010110100011010001,
    24'b000001100110100011001101,
    24'b000111110101000010000101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111101001110000111010110,
    24'b111100101110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110001011011000,
    24'b111011111110000111010110,
    24'b111100001110000111010111,
    24'b110110111101010011001110,
    24'b000000000000000000000000,
    24'b000000000000110100110101,
    24'b000100000110010010111010,
    24'b000000000110011111010011,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111010010,
    24'b000000000110011111001111,
    24'b000000010110011111001100,
    24'b000000010110010011001001,
    24'b000111010101100110011011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111011111110001111011000,
    24'b111100101110001011010011,
    24'b111100001110001011010111,
    24'b111100001110001011011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100101110000111011000,
    24'b111011101110000011010111,
    24'b101010011010000010100000,
    24'b000000000000000000000000,
    24'b000000000001001101000100,
    24'b000010010110001011000100,
    24'b000000000110011111001011,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011111010001,
    24'b000000000110011111001111,
    24'b000000100110011111001101,
    24'b000000010110010111001100,
    24'b000111010101111010101011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111011001101111111011000,
    24'b111100011110000111010111,
    24'b111100001110001011011001,
    24'b111100001110001011011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100001101111111010111,
    24'b111011111110000011011001,
    24'b001111110011010100110101,
    24'b000000000000000000000000,
    24'b000011010010111101100010,
    24'b000010010110001111000111,
    24'b000000000110011111001100,
    24'b000000010110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000100110011111001110,
    24'b000000110110011011001111,
    24'b000101100101111110110101,
    24'b000000000000111000101110,
    24'b000000000000000000000000,
    24'b101111011011001010101000,
    24'b111011111110000011011010,
    24'b111100001110000111011001,
    24'b111100001110001011011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100111110001011011010,
    24'b111011101110000111011001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000111110100111010001000,
    24'b000010010110010011001001,
    24'b000000010110011011010010,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100011001110,
    24'b000000000110011111001110,
    24'b000000100110011111001111,
    24'b000000100110010011001111,
    24'b000100000110001110111110,
    24'b000000100001111001001000,
    24'b000000000000000000000000,
    24'b011100110110100101100001,
    24'b111011111110001011011010,
    24'b111100101110010011011011,
    24'b111011111110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000011010111,
    24'b111011111101111011010110,
    24'b111001011101011111010010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000110110101101110100011,
    24'b000001100110011111001100,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110100011001100,
    24'b000000000110011111001101,
    24'b000000010110011011010000,
    24'b000001010110100011010010,
    24'b000001110110011011000110,
    24'b000101010100101110000111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111011101110011011011101,
    24'b111011111110000111011000,
    24'b111100001110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000011011000,
    24'b111100111110001011011010,
    24'b101101111010110010100110,
    24'b000000000000000000000000,
    24'b000000000000110000111000,
    24'b000110000110010011000000,
    24'b000001000110100011010000,
    24'b000000010110011011001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110100011001100,
    24'b000000000110011011001101,
    24'b000000000110010111001111,
    24'b000001100110100111010011,
    24'b000000010110011011001110,
    24'b001000010110001010101110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b110011111100100011000010,
    24'b111011111110001011011001,
    24'b111100101110001111011010,
    24'b111100011110000011010110,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110001011011001,
    24'b111100101110000111011000,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011011010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000011110010100101100010,
    24'b000011100110001111001010,
    24'b000000010110101011010101,
    24'b000000000110100011001101,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000001100110100111010000,
    24'b000000010110011111010101,
    24'b000101010110011011001001,
    24'b000001000001111001001011,
    24'b000000000000000000000000,
    24'b011000010101100001010111,
    24'b111010111101111011010101,
    24'b111100011110001111011001,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111011000,
    24'b111100111110000111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111011101110001111010110,
    24'b111100101110000011011001,
    24'b111101011110000011011000,
    24'b111100001110001011010110,
    24'b110111011101001011001100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000110100101001010011111,
    24'b000010000110001111001110,
    24'b000000010110011111010110,
    24'b000000110110011111010001,
    24'b000000010110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000100110011111010001,
    24'b000000010110100011010011,
    24'b000000010110011011010100,
    24'b000010110110010011001000,
    24'b000101010100101010001010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111011111110001111011101,
    24'b111100001110000111011000,
    24'b111100111110001111010110,
    24'b111100111110000111010101,
    24'b111100101110000111010110,
    24'b111100001110001011010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110001011010011,
    24'b111100111110001011010001,
    24'b111100011110000111010110,
    24'b111011101110010011100000,
    24'b011011000110100001100100,
    24'b000000000000000000000000,
    24'b000000000001011100111110,
    24'b000110000110101011000001,
    24'b000001000110001011000111,
    24'b000000000110011111010011,
    24'b000000010110011011010001,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000100110011111010001,
    24'b000000100110100011010010,
    24'b000000000110011011010011,
    24'b000001010110010111010000,
    24'b000001110110001111001000,
    24'b000110000110001110110101,
    24'b000000100001001100110100,
    24'b000000000000000000000000,
    24'b011110010110111001101001,
    24'b111011111110001011011010,
    24'b111100011110000011010110,
    24'b111100101110001011010011,
    24'b111100011110001011010101,
    24'b111100001110001011010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111101001101111111011001,
    24'b111100011110000111010010,
    24'b111011111110000111010111,
    24'b111010001101101111011100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000100000100100110001100,
    24'b000000000110100111001011,
    24'b000000110110010111000101,
    24'b000000010110100011010000,
    24'b000000010110011011010001,
    24'b000000010110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010011,
    24'b000001110110011011010000,
    24'b000001110110010111001010,
    24'b000011000110010011000101,
    24'b000011000011110001110110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111011001110001111011110,
    24'b111011001101111111010011,
    24'b111100001110001011010110,
    24'b111100011110000011010101,
    24'b111100111110001011011010,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101101111111011001,
    24'b111100011110010011011011,
    24'b111011101110000011011000,
    24'b011010000101011101010111,
    24'b000000000000000000000000,
    24'b000000010001000000101110,
    24'b000110010110010110111011,
    24'b000000000110110011011000,
    24'b000000110110011011001001,
    24'b000000000110100011001101,
    24'b000000000110011011010001,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000100110011011010011,
    24'b000000100110011011010110,
    24'b000000010110011011001110,
    24'b000001110110011011001111,
    24'b000110100110010010111100,
    24'b000000000001010100111100,
    24'b000000000000000000000000,
    24'b010001110100000100111110,
    24'b111010111110000111011000,
    24'b111100001110001011010101,
    24'b111100101110000011011000,
    24'b111100101101111111011001,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111001111,
    24'b111011101110000011011010,
    24'b111000101101001111001110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000101100100100010001010,
    24'b000010110110001111000010,
    24'b000000110110010011010100,
    24'b000000010110011011010000,
    24'b000000010110011011001101,
    24'b000000000110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110010111010111,
    24'b000000100110011111010110,
    24'b000000010110100111010011,
    24'b000011100110101111001000,
    24'b000101000100101110010100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101111111011010110110000,
    24'b111110001110011011011110,
    24'b111101011110001111011100,
    24'b111100001110001011010010,
    24'b111100111110000111010111,
    24'b111100011110000111011000,
    24'b111100111110001011011000,
    24'b111100111110000111010101,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110001011011000,
    24'b111011101101111111010011,
    24'b111100111110001011010110,
    24'b111100001101101111001000,
    24'b111011001110001111010100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000100001101001001010,
    24'b000101010110001110111101,
    24'b000001100110011011001100,
    24'b000000110110010111010010,
    24'b000000010110011011010001,
    24'b000000010110011011001111,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010001,
    24'b000000100110010111010100,
    24'b000000000110011111010010,
    24'b000001000110010111001000,
    24'b000110000110001011000001,
    24'b000010000010101001010110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111001011110000111011000,
    24'b111011001110010011010111,
    24'b111101011101111011010111,
    24'b111100111110000111010110,
    24'b111100001110001011011001,
    24'b111100011110000011010110,
    24'b111101001110000011010101,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100101110001011010101,
    24'b111011011101110111010000,
    24'b111011011101110111011000,
    24'b011010100110010101011111,
    24'b000000000000000000000000,
    24'b000000000000101000101000,
    24'b000110000101011010100000,
    24'b000001110110011111001011,
    24'b000001100110101111010101,
    24'b000000000110010111001111,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110011011001110,
    24'b000001000110010011010010,
    24'b000000000110001111001111,
    24'b000000110110100011010001,
    24'b000011010110011011001101,
    24'b000101110101110110110011,
    24'b000000000001001000110011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b111001001101111111010101,
    24'b111110011101110011011000,
    24'b111100011110000111011000,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100111110001011011010,
    24'b111100111110001011011000,
    24'b111100111110000111010111,
    24'b111100101110000111011000,
    24'b111101001110010011011011,
    24'b101100011010011110100101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000101100100000101111101,
    24'b000010100110011111001000,
    24'b000000000110011011010000,
    24'b000000100110011111010001,
    24'b000000100110011111010001,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000010110011011010011,
    24'b000000100110010111010100,
    24'b000000100110011011010011,
    24'b000000000110010111001101,
    24'b000001110110101011001110,
    24'b000010000110100011001001,
    24'b000101110101000010010101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010100010100011001000110,
    24'b111010111110001011011001,
    24'b111100101110010111011101,
    24'b111100111110000011010101,
    24'b111100101110000011010110,
    24'b111100001110000111011010,
    24'b111100011110000111010111,
    24'b111100101110000111010110,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001101111011010100,
    24'b111101001110001011011000,
    24'b111101001110001111011001,
    24'b111100011110001111011100,
    24'b110011101100001010111101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000001010010100101011100,
    24'b000101000110001010111001,
    24'b000000110110010111001100,
    24'b000000000110011111010100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010100,
    24'b000000000110011111010010,
    24'b000000000110011111010000,
    24'b000000010110011011001100,
    24'b000000110110011011001101,
    24'b000001000110100011000011,
    24'b000011110110010011001110,
    24'b000100110100001010001010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010101000101011101011001,
    24'b111010111101111111011001,
    24'b111101111110000011010101,
    24'b111110001110010011011011,
    24'b111011001110000111011101,
    24'b111011111110000111010110,
    24'b111100101110000111010100,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110001011011000,
    24'b111100111110001011011000,
    24'b111100011101111111010100,
    24'b111101011110001111010110,
    24'b111100011101111111010011,
    24'b111101001110010011011100,
    24'b110010001011111010111011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000100001110000111111,
    24'b000100100110001010110101,
    24'b000000110110011111001101,
    24'b000000110110011011001011,
    24'b000000010110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110101011001100,
    24'b000000000110100011001110,
    24'b000001010110010111010010,
    24'b000001100110001111010011,
    24'b000001010110001111010000,
    24'b000000100110100011010001,
    24'b000011000110001111000011,
    24'b000100010011110001110010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010011110100010101000001,
    24'b111100101101101111001111,
    24'b111101111110000111011010,
    24'b111011001110001011011111,
    24'b111100001110001011010111,
    24'b111100101110001011010100,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110000011010110,
    24'b111100001110000011010110,
    24'b111101001110001111010101,
    24'b111100011110000011010000,
    24'b111101111110011011011000,
    24'b101110101010110110100101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001011100111111,
    24'b000110010101110110101111,
    24'b000010000110010111001000,
    24'b000000100110101111010010,
    24'b000000000110100011010001,
    24'b000000000110010111001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000010110011111010101,
    24'b000000010110011111010101,
    24'b000000100110011111001110,
    24'b000001000110011011001011,
    24'b000001100110010111001111,
    24'b000011110110001111000100,
    24'b000100000011111101111100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001010000010001100100110,
    24'b111010001101111111011011,
    24'b111100011110000011010110,
    24'b111110001110010111010111,
    24'b111101001110000111010011,
    24'b111100101110000111010111,
    24'b111100001110001011011001,
    24'b111100001110001011010101,
    24'b111100101110001011010011,
    24'b111101011110000111011000,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110001011010101,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011001,
    24'b111100111110000011011001,
    24'b111100101110000111010110,
    24'b111100101110001011010101,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100101110000111011000,
    24'b111100101110000111011001,
    24'b111011111110000111011000,
    24'b111100111110001011010010,
    24'b111100101110001011010110,
    24'b111011011101111111011100,
    24'b111100011110001011011101,
    24'b111100001101110011011000,
    24'b111011101110001111010100,
    24'b100011001000011110000001,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000010001101100111110,
    24'b000010000110000010110100,
    24'b000001100110010011000001,
    24'b000000010110011011001011,
    24'b000000000110011011001110,
    24'b000000010110100011001110,
    24'b000000010110100011001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010000,
    24'b000000110110100011010100,
    24'b000000110110010111001101,
    24'b000000010110011011010000,
    24'b000001110110101111010100,
    24'b000100110110000110111011,
    24'b000101000100011110001010,
    24'b000000000000101000101000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b101011101010100010101000,
    24'b111010011101111111011010,
    24'b111011111101110111010011,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000111010100,
    24'b111100101110001011010101,
    24'b111100101110000011010110,
    24'b111100001110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100101110000111010111,
    24'b111100111110000111010110,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100011110000111011001,
    24'b111100001110001011010111,
    24'b111100001110001011010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000011011000,
    24'b111101111101111011011010,
    24'b111101111101111111010100,
    24'b111101001110000111010101,
    24'b111100111110000011011001,
    24'b111100001110000011010001,
    24'b111011101101101111010010,
    24'b010000110011110000110110,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000110001111101000100,
    24'b000100100110001110110011,
    24'b000010010110011011000111,
    24'b000001110110100011001111,
    24'b000000000110010111010001,
    24'b000000000110100011010110,
    24'b000000000110011011010011,
    24'b000000010110011011010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000010110100011001111,
    24'b000000000110011111001100,
    24'b000000010110100011010101,
    24'b000000110110100011010001,
    24'b000000000110011011001101,
    24'b000000000110011111010001,
    24'b000001000110010111010001,
    24'b000011100110010111001001,
    24'b000101010101001010010111,
    24'b000000000001010100111000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010100000100011000111110,
    24'b111001011101011111010000,
    24'b111100001110000111011010,
    24'b111011111101111011010100,
    24'b111101011110010011011010,
    24'b111100101110000111011000,
    24'b111100111110010011010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100111110000111010111,
    24'b111101001110000011010111,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100001110001011010111,
    24'b111100001110001011011001,
    24'b111100001110001011011001,
    24'b111100001110001011011001,
    24'b111100001110001011010111,
    24'b111100111110000111010111,
    24'b111100111110000011010111,
    24'b111010101110010111010101,
    24'b111011111110010011011010,
    24'b111100111110000011011101,
    24'b111100111110001011100011,
    24'b100111001001010110010101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000010010011010101101010,
    24'b000101110110010110110110,
    24'b000001000110101011010000,
    24'b000000100110011011010000,
    24'b000000010110011011010010,
    24'b000000000110011111010101,
    24'b000000010110101011011000,
    24'b000000000110010111010011,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001110,
    24'b000000000110011111001101,
    24'b000000000110100011010010,
    24'b000000000110100011010000,
    24'b000000000110100011001011,
    24'b000000010110100011001010,
    24'b000000100110011011001101,
    24'b000000100110011011001110,
    24'b000001100110011011000110,
    24'b000110110110001010101101,
    24'b000010100010101101010100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b011011000110010001100100,
    24'b111000111101100011010001,
    24'b111011111110000011011100,
    24'b111011111110000011011100,
    24'b111011011110000111010101,
    24'b111101111110001111011010,
    24'b111101001110000011010111,
    24'b111101001110000011010111,
    24'b111101001110000011010111,
    24'b111100111101111111010110,
    24'b111100111110000011010111,
    24'b111100111110000111011000,
    24'b111100111110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111010111,
    24'b111100101110000111011000,
    24'b111100101110001111011001,
    24'b111011111110001011011001,
    24'b111011111110000111011000,
    24'b111011111101111011010101,
    24'b111100101101111111011001,
    24'b111100101110000111011011,
    24'b111010011110010111011011,
    24'b101011001010101110011110,
    24'b001011110010011000011111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001010000111000,
    24'b000011010101000010010111,
    24'b000001110110011111000001,
    24'b000000000110010111001100,
    24'b000000110110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000000110011011010001,
    24'b000000000110011011001111,
    24'b000000000110011111010000,
    24'b000000000110011011010000,
    24'b000000110110011011001101,
    24'b000000010110011111001100,
    24'b000000000110011111001110,
    24'b000000000110010111001110,
    24'b000010000110011011001010,
    24'b000101010110010010111011,
    24'b000110010100111110010010,
    24'b000000000001011001000100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010101110100101101001101,
    24'b110001011011100110111001,
    24'b111011001110010011011001,
    24'b111101011110011011011100,
    24'b111011101101111111010100,
    24'b111100011110001011010111,
    24'b111100011110001011010111,
    24'b111100011110000111010111,
    24'b111100011110000111010111,
    24'b111100001110001011011001,
    24'b111100101110000111011001,
    24'b111100111110000111010111,
    24'b111100111110000111010111,
    24'b111100111110000111010101,
    24'b111100111110000011010100,
    24'b111100101110000111010101,
    24'b111011111110001111011010,
    24'b111011001110001011011000,
    24'b111011001101111011011000,
    24'b111001011101001011010000,
    24'b100101101000000110000101,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000001100011000101011110,
    24'b000111000110000110110010,
    24'b000010000110011011001011,
    24'b000000100110100111001010,
    24'b000000100110011111010000,
    24'b000000010110100011010001,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001101,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011011010011,
    24'b000000100110011011001110,
    24'b000000010110011011010010,
    24'b000000000110011011010100,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000100110010011001101,
    24'b000001010110011011010000,
    24'b000000100110010111010110,
    24'b000001010110010011001111,
    24'b000110100110001110111010,
    24'b000110000011111001111101,
    24'b000000010001001000110111,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b010110010101011101010000,
    24'b101011001010011110011111,
    24'b110110111101001111001010,
    24'b111001111101111111010101,
    24'b111011001110010111011011,
    24'b111011001110010011011011,
    24'b111100001110000111011010,
    24'b111100001110000111011011,
    24'b111100011110000111011011,
    24'b111100011110000111011001,
    24'b111100011110001011011000,
    24'b111100011110000111010101,
    24'b111001001101011011001100,
    24'b110011011100010010111011,
    24'b011111000111010001101110,
    24'b001100010010101100101010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000100000101100,
    24'b000001110010001101011011,
    24'b000110010101101110101000,
    24'b000000110110001111000001,
    24'b000010010110011111010001,
    24'b000010000110001111001001,
    24'b000001010110100011001010,
    24'b000000000110011011010010,
    24'b000000000110011111001110,
    24'b000000000110011011010001,
    24'b000000010110011011010000,
    24'b000000010110011011001110,
    24'b000000000110011111001111,
    24'b000000000110011011010001,
    24'b000000000110011111010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110100011010001,
    24'b000000000110011111001111,
    24'b000000000110011111001101,
    24'b000000010110011011010000,
    24'b000000100110011011010010,
    24'b000001000110010111001110,
    24'b000001010110011111001010,
    24'b000001110110010111000101,
    24'b000110110110100011000000,
    24'b000101110100101010001100,
    24'b000001010001111101001011,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b001101010011000100101101,
    24'b010000110011111100111110,
    24'b010001110100010001000011,
    24'b010001010100001101000011,
    24'b001110110011110000111010,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000001010100110110,
    24'b000010110011100001101111,
    24'b000110010101101010101010,
    24'b000100010110010111000101,
    24'b000001000110000111001000,
    24'b000000110110010011001011,
    24'b000001010110011011010000,
    24'b000001100110100011010110,
    24'b000000110110011111010110,
    24'b000000010110100011010001,
    24'b000000000110011111001100,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001110,
    24'b000000000110011111001101,
    24'b000000000110011111010000,
    24'b000000010110011011010010,
    24'b000001000110011011010011,
    24'b000001000110011111001111,
    24'b000000000110110011001110,
    24'b000000010110110011001111,
    24'b000010110110011111001110,
    24'b000101110110001011000001,
    24'b000111110101111010101011,
    24'b000011100100100010000010,
    24'b000010100010100001010011,
    24'b000000000000111100110100,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000000000000000,
    24'b000000000000101100101011,
    24'b000000000001110001000111,
    24'b000010100011010101101110,
    24'b000110010101001010011001,
    24'b000100000110010111000010,
    24'b000011100110100011001001,
    24'b000010000110101011001110,
    24'b000000000110010011001001,
    24'b000000000110100011001100,
    24'b000000010110011011001110,
    24'b000000110110010111010000,
    24'b000000100110011011010011,
    24'b000000110110011111010110,
    24'b000000010110011111010010,
    24'b000000000110011111001110,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110100011001110,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010011,
    24'b000000000110011011010010,
    24'b000000010110011011010010,
    24'b000000000110011111001110,
    24'b000000000110100111001011,
    24'b000000000110100111001100,
    24'b000000000110010111010001,
    24'b000001000110010011010101,
    24'b000001110110010111000110,
    24'b000011010110001010111100,
    24'b000100110101110110101011,
    24'b000101100101011010011001,
    24'b000100000100011110000010,
    24'b000100000011111101111010,
    24'b000011110011100101110111,
    24'b000011100011100001101111,
    24'b000011110011100101101101,
    24'b000100000011110001110011,
    24'b000101100100001110000001,
    24'b000101010101000010011011,
    24'b000101100101100110101010,
    24'b000100110101111010110100,
    24'b000011010110001010111010,
    24'b000010000110010111000011,
    24'b000001010110010111001101,
    24'b000000110110010111001111,
    24'b000000110110011011001101,
    24'b000000010110011111001011,
    24'b000000110110011011001011,
    24'b000000110110011011001010,
    24'b000000110110011011001101,
    24'b000000010110010111010000,
    24'b000000010110011011010001,
    24'b000000010110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011011010010,
    24'b000000010110010111010100,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000000110011111001111,
    24'b000000010110011011001101,
    24'b000000110110011011001011,
    24'b000000100110011011001011,
    24'b000000010110011011001010,
    24'b000000010110011011001001,
    24'b000000100110011111001010,
    24'b000001000110100111001101,
    24'b000001100110100111001011,
    24'b000001110110100011000110,
    24'b000001110110011111000011,
    24'b000001100110011011000001,
    24'b000001110110011111000100,
    24'b000001010110011011000101,
    24'b000001000110010011001000,
    24'b000001000110011011001110,
    24'b000000110110011111010000,
    24'b000000010110100111001101,
    24'b000000000110100011001101,
    24'b000000000110011111010001,
    24'b000000000110011111001110,
    24'b000000000110011111001110,
    24'b000000000110011111010001,
    24'b000000000110011011010011,
    24'b000000000110011011010100,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000010110011011010000,
    24'b000000010110011011001111,
    24'b000000010110011111001111,
    24'b000000010110011111010000,
    24'b000000010110011011010001,
    24'b000000100110011011010010,
    24'b000000010110011011010011,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110100011001101,
    24'b000000010110011111001111,
    24'b000000010110011111010000,
    24'b000000000110010111010000,
    24'b000000100110011111010001,
    24'b000000110110011011010001,
    24'b000000110110011111001110,
    24'b000000110110100011001110,
    24'b000001010110011111001111,
    24'b000001010110011011010000,
    24'b000000110110010111001101,
    24'b000000100110011111001100,
    24'b000000110110011011001111,
    24'b000000110110011111010011,
    24'b000000010110100011010101,
    24'b000000000110100011001111,
    24'b000000010110011111001110,
    24'b000000100110010111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010010,
    24'b000000010110011011010011,
    24'b000000010110011111010010,
    24'b000000010110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011011010001,
    24'b000000000110011111010001,
    24'b000000000110011011010011,
    24'b000000000110011011010010,
    24'b000000010110011011010011,
    24'b000000100110011111010100,
    24'b000000100110011011010011,
    24'b000000110110010111010010,
    24'b000001000110010111010000,
    24'b000001010110010111010010,
    24'b000000100110010111010010,
    24'b000000010110011011010011,
    24'b000000010110010111010011,
    24'b000000000110010111010000,
    24'b000000000110011111001101,
    24'b000000000110011111001011,
    24'b000000010110011011001110,
    24'b000000010110011011010001,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011010000,
    24'b000000000110011111001110,
    24'b000000000110011111001111,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111001111,
    24'b000000000110011111001111,
    24'b000000000110011011010001,
    24'b000000000110011011010001,
    24'b000000010110011111010011,
    24'b000000010110011011010010,
    24'b000000010110011011010010,
    24'b000000100110010111010000,
    24'b000000100110010111010000,
    24'b000000000110011011010010,
    24'b000000000110011111010100,
    24'b000000010110011011010010,
    24'b000000010110011011001111,
    24'b000000010110011111001100,
    24'b000000000110100011001011,
    24'b000000000110011111001111,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000010110011011001110,
    24'b000000000110011111001100,
    24'b000000000110011111001101,
    24'b000000010110100011001111,
    24'b000000100110100111010010,
    24'b000000000110100111010010,
    24'b000000000110100011010011,
    24'b000000010110100011010001,
    24'b000000000110011111010000,
    24'b000000010110100111010100,
    24'b000000000110100111010110,
    24'b000000010110011111010011,
    24'b000000000110011111010000,
    24'b000000010110100011001111,
    24'b000000010110100011001111,
    24'b000000000110011111010000,
    24'b000000000110011011010010,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000,
    24'b000000000110011111010000
};


assign mem = memory;

endmodule
