library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity sumador_1bit is
    Port ( A    : in  STD_LOGIC;
           B    : in  STD_LOGIC;
           Cin  : in  STD_LOGIC;
           S    : out STD_LOGIC;
           Cout : out STD_LOGIC);
end sumador_1bit;

architecture Behavioral of sumador_1bit is
begin
    S    <= A XOR B XOR Cin;
    Cout <= (A AND B) OR (A AND Cin) OR (B AND Cin);
end Behavioral;